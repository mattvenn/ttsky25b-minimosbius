VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mosbius
  CLASS BLOCK ;
  FOREIGN tt_um_mosbius ;
  ORIGIN 0.000 0.000 ;
  SIZE 493.120 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.330 9.400 2.530 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.190 9.400 21.390 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.050 9.400 40.250 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.910 9.400 59.110 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.770 9.400 77.970 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.630 9.400 96.830 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.490 9.400 115.690 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 133.350 9.400 134.550 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.210 9.400 153.410 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.070 9.400 172.270 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.930 9.400 191.130 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.790 9.400 209.990 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.650 9.400 228.850 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.510 9.400 247.710 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 265.370 9.400 266.570 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.230 9.400 285.430 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 303.090 9.400 304.290 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.950 9.400 323.150 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 340.810 9.400 342.010 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.670 9.400 360.870 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.530 9.400 379.730 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 397.390 9.400 398.590 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.250 9.400 417.450 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 435.110 9.400 436.310 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 453.970 9.400 455.170 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 472.830 9.400 474.030 220.970 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2.930 9.400 4.130 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.790 9.400 22.990 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.650 9.400 41.850 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.510 9.400 60.710 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.370 9.400 79.570 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.230 9.400 98.430 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.090 9.400 117.290 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.950 9.400 136.150 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.810 9.400 155.010 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 172.670 9.400 173.870 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.530 9.400 192.730 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 210.390 9.400 211.590 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 229.250 9.400 230.450 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.110 9.400 249.310 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 266.970 9.400 268.170 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 285.830 9.400 287.030 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.690 9.400 305.890 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.550 9.400 324.750 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 342.410 9.400 343.610 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 361.270 9.400 362.470 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 380.130 9.400 381.330 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 398.990 9.400 400.190 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 417.850 9.400 419.050 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.710 9.400 437.910 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 455.570 9.400 456.770 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.430 9.400 475.630 220.970 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.530 9.400 5.730 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.390 9.400 24.590 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.250 9.400 43.450 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.110 9.400 62.310 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.970 9.400 81.170 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.830 9.400 100.030 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.690 9.400 118.890 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.550 9.400 137.750 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 155.410 9.400 156.610 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.270 9.400 175.470 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 193.130 9.400 194.330 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.990 9.400 213.190 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 230.850 9.400 232.050 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.710 9.400 250.910 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.570 9.400 269.770 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 287.430 9.400 288.630 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 306.290 9.400 307.490 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.150 9.400 326.350 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.010 9.400 345.210 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 362.870 9.400 364.070 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.730 9.400 382.930 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.590 9.400 401.790 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 419.450 9.400 420.650 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 438.310 9.400 439.510 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 457.170 9.400 458.370 220.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.030 9.400 477.230 220.970 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 0.500 219.395 3.640 221.000 ;
        RECT 0.500 219.390 3.180 219.395 ;
        RECT 0.500 213.955 491.700 216.785 ;
        RECT 0.500 208.515 491.700 211.345 ;
        RECT 0.500 204.300 491.700 205.905 ;
      LAYER li1 ;
        RECT 0.680 0.820 491.510 223.615 ;
      LAYER met1 ;
        RECT 0.690 0.000 491.510 225.750 ;
      LAYER met2 ;
        RECT 1.200 0.000 490.940 225.750 ;
      LAYER met3 ;
        RECT 0.850 0.000 491.320 225.750 ;
      LAYER met4 ;
        RECT 6.410 224.360 14.630 225.750 ;
        RECT 15.730 224.360 17.390 225.750 ;
        RECT 18.490 224.360 20.150 225.750 ;
        RECT 21.250 224.360 22.910 225.750 ;
        RECT 24.010 224.360 25.670 225.750 ;
        RECT 26.770 224.360 28.430 225.750 ;
        RECT 29.530 224.360 31.190 225.750 ;
        RECT 32.290 224.360 33.950 225.750 ;
        RECT 35.050 224.360 36.710 225.750 ;
        RECT 37.810 224.360 39.470 225.750 ;
        RECT 40.570 224.360 42.230 225.750 ;
        RECT 43.330 224.360 44.990 225.750 ;
        RECT 46.090 224.360 47.750 225.750 ;
        RECT 48.850 224.360 50.510 225.750 ;
        RECT 51.610 224.360 53.270 225.750 ;
        RECT 54.370 224.360 56.030 225.750 ;
        RECT 57.130 224.360 58.790 225.750 ;
        RECT 59.890 224.360 61.550 225.750 ;
        RECT 62.650 224.360 64.310 225.750 ;
        RECT 65.410 224.360 67.070 225.750 ;
        RECT 68.170 224.360 69.830 225.750 ;
        RECT 70.930 224.360 72.590 225.750 ;
        RECT 73.690 224.360 75.350 225.750 ;
        RECT 76.450 224.360 78.110 225.750 ;
        RECT 79.210 224.360 80.870 225.750 ;
        RECT 81.970 224.360 83.630 225.750 ;
        RECT 84.730 224.360 86.390 225.750 ;
        RECT 87.490 224.360 89.150 225.750 ;
        RECT 90.250 224.360 91.910 225.750 ;
        RECT 93.010 224.360 94.670 225.750 ;
        RECT 95.770 224.360 97.430 225.750 ;
        RECT 98.530 224.360 100.190 225.750 ;
        RECT 101.290 224.360 102.950 225.750 ;
        RECT 104.050 224.360 105.710 225.750 ;
        RECT 106.810 224.360 108.470 225.750 ;
        RECT 109.570 224.360 111.230 225.750 ;
        RECT 112.330 224.360 113.990 225.750 ;
        RECT 115.090 224.360 116.750 225.750 ;
        RECT 117.850 224.360 119.510 225.750 ;
        RECT 120.610 224.360 122.270 225.750 ;
        RECT 123.370 224.360 125.030 225.750 ;
        RECT 126.130 224.360 127.790 225.750 ;
        RECT 128.890 224.360 130.550 225.750 ;
        RECT 131.650 224.360 490.800 225.750 ;
        RECT 6.410 221.370 490.800 224.360 ;
        RECT 6.410 9.000 19.790 221.370 ;
        RECT 24.990 9.000 38.650 221.370 ;
        RECT 43.850 9.000 57.510 221.370 ;
        RECT 62.710 9.000 76.370 221.370 ;
        RECT 81.570 9.000 95.230 221.370 ;
        RECT 100.430 9.000 114.090 221.370 ;
        RECT 119.290 9.000 132.950 221.370 ;
        RECT 138.150 9.000 151.810 221.370 ;
        RECT 157.010 9.000 170.670 221.370 ;
        RECT 175.870 9.000 189.530 221.370 ;
        RECT 194.730 9.000 208.390 221.370 ;
        RECT 213.590 9.000 227.250 221.370 ;
        RECT 232.450 9.000 246.110 221.370 ;
        RECT 251.310 9.000 264.970 221.370 ;
        RECT 270.170 9.000 283.830 221.370 ;
        RECT 289.030 9.000 302.690 221.370 ;
        RECT 307.890 9.000 321.550 221.370 ;
        RECT 326.750 9.000 340.410 221.370 ;
        RECT 345.610 9.000 359.270 221.370 ;
        RECT 364.470 9.000 378.130 221.370 ;
        RECT 383.330 9.000 396.990 221.370 ;
        RECT 402.190 9.000 415.850 221.370 ;
        RECT 421.050 9.000 434.710 221.370 ;
        RECT 439.910 9.000 453.570 221.370 ;
        RECT 458.770 9.000 472.430 221.370 ;
        RECT 477.630 9.000 490.800 221.370 ;
        RECT 6.410 1.400 490.800 9.000 ;
        RECT 6.410 0.000 19.850 1.400 ;
        RECT 21.550 0.000 39.170 1.400 ;
        RECT 40.870 0.000 58.490 1.400 ;
        RECT 60.190 0.000 77.810 1.400 ;
        RECT 79.510 0.000 97.130 1.400 ;
        RECT 98.830 0.000 116.450 1.400 ;
        RECT 118.150 0.000 135.770 1.400 ;
        RECT 137.470 0.000 490.800 1.400 ;
  END
END tt_um_mosbius
END LIBRARY


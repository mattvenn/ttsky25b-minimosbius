magic
tech sky130A
magscale 1 2
timestamp 1757785414
<< pwell >>
rect -3811 -1367 3811 1367
<< mvnmos >>
rect -3583 109 -3383 1109
rect -3325 109 -3125 1109
rect -3067 109 -2867 1109
rect -2809 109 -2609 1109
rect -2551 109 -2351 1109
rect -2293 109 -2093 1109
rect -2035 109 -1835 1109
rect -1777 109 -1577 1109
rect -1519 109 -1319 1109
rect -1261 109 -1061 1109
rect -1003 109 -803 1109
rect -745 109 -545 1109
rect -487 109 -287 1109
rect -229 109 -29 1109
rect 29 109 229 1109
rect 287 109 487 1109
rect 545 109 745 1109
rect 803 109 1003 1109
rect 1061 109 1261 1109
rect 1319 109 1519 1109
rect 1577 109 1777 1109
rect 1835 109 2035 1109
rect 2093 109 2293 1109
rect 2351 109 2551 1109
rect 2609 109 2809 1109
rect 2867 109 3067 1109
rect 3125 109 3325 1109
rect 3383 109 3583 1109
rect -3583 -1109 -3383 -109
rect -3325 -1109 -3125 -109
rect -3067 -1109 -2867 -109
rect -2809 -1109 -2609 -109
rect -2551 -1109 -2351 -109
rect -2293 -1109 -2093 -109
rect -2035 -1109 -1835 -109
rect -1777 -1109 -1577 -109
rect -1519 -1109 -1319 -109
rect -1261 -1109 -1061 -109
rect -1003 -1109 -803 -109
rect -745 -1109 -545 -109
rect -487 -1109 -287 -109
rect -229 -1109 -29 -109
rect 29 -1109 229 -109
rect 287 -1109 487 -109
rect 545 -1109 745 -109
rect 803 -1109 1003 -109
rect 1061 -1109 1261 -109
rect 1319 -1109 1519 -109
rect 1577 -1109 1777 -109
rect 1835 -1109 2035 -109
rect 2093 -1109 2293 -109
rect 2351 -1109 2551 -109
rect 2609 -1109 2809 -109
rect 2867 -1109 3067 -109
rect 3125 -1109 3325 -109
rect 3383 -1109 3583 -109
<< mvndiff >>
rect -3641 1097 -3583 1109
rect -3641 121 -3629 1097
rect -3595 121 -3583 1097
rect -3641 109 -3583 121
rect -3383 1097 -3325 1109
rect -3383 121 -3371 1097
rect -3337 121 -3325 1097
rect -3383 109 -3325 121
rect -3125 1097 -3067 1109
rect -3125 121 -3113 1097
rect -3079 121 -3067 1097
rect -3125 109 -3067 121
rect -2867 1097 -2809 1109
rect -2867 121 -2855 1097
rect -2821 121 -2809 1097
rect -2867 109 -2809 121
rect -2609 1097 -2551 1109
rect -2609 121 -2597 1097
rect -2563 121 -2551 1097
rect -2609 109 -2551 121
rect -2351 1097 -2293 1109
rect -2351 121 -2339 1097
rect -2305 121 -2293 1097
rect -2351 109 -2293 121
rect -2093 1097 -2035 1109
rect -2093 121 -2081 1097
rect -2047 121 -2035 1097
rect -2093 109 -2035 121
rect -1835 1097 -1777 1109
rect -1835 121 -1823 1097
rect -1789 121 -1777 1097
rect -1835 109 -1777 121
rect -1577 1097 -1519 1109
rect -1577 121 -1565 1097
rect -1531 121 -1519 1097
rect -1577 109 -1519 121
rect -1319 1097 -1261 1109
rect -1319 121 -1307 1097
rect -1273 121 -1261 1097
rect -1319 109 -1261 121
rect -1061 1097 -1003 1109
rect -1061 121 -1049 1097
rect -1015 121 -1003 1097
rect -1061 109 -1003 121
rect -803 1097 -745 1109
rect -803 121 -791 1097
rect -757 121 -745 1097
rect -803 109 -745 121
rect -545 1097 -487 1109
rect -545 121 -533 1097
rect -499 121 -487 1097
rect -545 109 -487 121
rect -287 1097 -229 1109
rect -287 121 -275 1097
rect -241 121 -229 1097
rect -287 109 -229 121
rect -29 1097 29 1109
rect -29 121 -17 1097
rect 17 121 29 1097
rect -29 109 29 121
rect 229 1097 287 1109
rect 229 121 241 1097
rect 275 121 287 1097
rect 229 109 287 121
rect 487 1097 545 1109
rect 487 121 499 1097
rect 533 121 545 1097
rect 487 109 545 121
rect 745 1097 803 1109
rect 745 121 757 1097
rect 791 121 803 1097
rect 745 109 803 121
rect 1003 1097 1061 1109
rect 1003 121 1015 1097
rect 1049 121 1061 1097
rect 1003 109 1061 121
rect 1261 1097 1319 1109
rect 1261 121 1273 1097
rect 1307 121 1319 1097
rect 1261 109 1319 121
rect 1519 1097 1577 1109
rect 1519 121 1531 1097
rect 1565 121 1577 1097
rect 1519 109 1577 121
rect 1777 1097 1835 1109
rect 1777 121 1789 1097
rect 1823 121 1835 1097
rect 1777 109 1835 121
rect 2035 1097 2093 1109
rect 2035 121 2047 1097
rect 2081 121 2093 1097
rect 2035 109 2093 121
rect 2293 1097 2351 1109
rect 2293 121 2305 1097
rect 2339 121 2351 1097
rect 2293 109 2351 121
rect 2551 1097 2609 1109
rect 2551 121 2563 1097
rect 2597 121 2609 1097
rect 2551 109 2609 121
rect 2809 1097 2867 1109
rect 2809 121 2821 1097
rect 2855 121 2867 1097
rect 2809 109 2867 121
rect 3067 1097 3125 1109
rect 3067 121 3079 1097
rect 3113 121 3125 1097
rect 3067 109 3125 121
rect 3325 1097 3383 1109
rect 3325 121 3337 1097
rect 3371 121 3383 1097
rect 3325 109 3383 121
rect 3583 1097 3641 1109
rect 3583 121 3595 1097
rect 3629 121 3641 1097
rect 3583 109 3641 121
rect -3641 -121 -3583 -109
rect -3641 -1097 -3629 -121
rect -3595 -1097 -3583 -121
rect -3641 -1109 -3583 -1097
rect -3383 -121 -3325 -109
rect -3383 -1097 -3371 -121
rect -3337 -1097 -3325 -121
rect -3383 -1109 -3325 -1097
rect -3125 -121 -3067 -109
rect -3125 -1097 -3113 -121
rect -3079 -1097 -3067 -121
rect -3125 -1109 -3067 -1097
rect -2867 -121 -2809 -109
rect -2867 -1097 -2855 -121
rect -2821 -1097 -2809 -121
rect -2867 -1109 -2809 -1097
rect -2609 -121 -2551 -109
rect -2609 -1097 -2597 -121
rect -2563 -1097 -2551 -121
rect -2609 -1109 -2551 -1097
rect -2351 -121 -2293 -109
rect -2351 -1097 -2339 -121
rect -2305 -1097 -2293 -121
rect -2351 -1109 -2293 -1097
rect -2093 -121 -2035 -109
rect -2093 -1097 -2081 -121
rect -2047 -1097 -2035 -121
rect -2093 -1109 -2035 -1097
rect -1835 -121 -1777 -109
rect -1835 -1097 -1823 -121
rect -1789 -1097 -1777 -121
rect -1835 -1109 -1777 -1097
rect -1577 -121 -1519 -109
rect -1577 -1097 -1565 -121
rect -1531 -1097 -1519 -121
rect -1577 -1109 -1519 -1097
rect -1319 -121 -1261 -109
rect -1319 -1097 -1307 -121
rect -1273 -1097 -1261 -121
rect -1319 -1109 -1261 -1097
rect -1061 -121 -1003 -109
rect -1061 -1097 -1049 -121
rect -1015 -1097 -1003 -121
rect -1061 -1109 -1003 -1097
rect -803 -121 -745 -109
rect -803 -1097 -791 -121
rect -757 -1097 -745 -121
rect -803 -1109 -745 -1097
rect -545 -121 -487 -109
rect -545 -1097 -533 -121
rect -499 -1097 -487 -121
rect -545 -1109 -487 -1097
rect -287 -121 -229 -109
rect -287 -1097 -275 -121
rect -241 -1097 -229 -121
rect -287 -1109 -229 -1097
rect -29 -121 29 -109
rect -29 -1097 -17 -121
rect 17 -1097 29 -121
rect -29 -1109 29 -1097
rect 229 -121 287 -109
rect 229 -1097 241 -121
rect 275 -1097 287 -121
rect 229 -1109 287 -1097
rect 487 -121 545 -109
rect 487 -1097 499 -121
rect 533 -1097 545 -121
rect 487 -1109 545 -1097
rect 745 -121 803 -109
rect 745 -1097 757 -121
rect 791 -1097 803 -121
rect 745 -1109 803 -1097
rect 1003 -121 1061 -109
rect 1003 -1097 1015 -121
rect 1049 -1097 1061 -121
rect 1003 -1109 1061 -1097
rect 1261 -121 1319 -109
rect 1261 -1097 1273 -121
rect 1307 -1097 1319 -121
rect 1261 -1109 1319 -1097
rect 1519 -121 1577 -109
rect 1519 -1097 1531 -121
rect 1565 -1097 1577 -121
rect 1519 -1109 1577 -1097
rect 1777 -121 1835 -109
rect 1777 -1097 1789 -121
rect 1823 -1097 1835 -121
rect 1777 -1109 1835 -1097
rect 2035 -121 2093 -109
rect 2035 -1097 2047 -121
rect 2081 -1097 2093 -121
rect 2035 -1109 2093 -1097
rect 2293 -121 2351 -109
rect 2293 -1097 2305 -121
rect 2339 -1097 2351 -121
rect 2293 -1109 2351 -1097
rect 2551 -121 2609 -109
rect 2551 -1097 2563 -121
rect 2597 -1097 2609 -121
rect 2551 -1109 2609 -1097
rect 2809 -121 2867 -109
rect 2809 -1097 2821 -121
rect 2855 -1097 2867 -121
rect 2809 -1109 2867 -1097
rect 3067 -121 3125 -109
rect 3067 -1097 3079 -121
rect 3113 -1097 3125 -121
rect 3067 -1109 3125 -1097
rect 3325 -121 3383 -109
rect 3325 -1097 3337 -121
rect 3371 -1097 3383 -121
rect 3325 -1109 3383 -1097
rect 3583 -121 3641 -109
rect 3583 -1097 3595 -121
rect 3629 -1097 3641 -121
rect 3583 -1109 3641 -1097
<< mvndiffc >>
rect -3629 121 -3595 1097
rect -3371 121 -3337 1097
rect -3113 121 -3079 1097
rect -2855 121 -2821 1097
rect -2597 121 -2563 1097
rect -2339 121 -2305 1097
rect -2081 121 -2047 1097
rect -1823 121 -1789 1097
rect -1565 121 -1531 1097
rect -1307 121 -1273 1097
rect -1049 121 -1015 1097
rect -791 121 -757 1097
rect -533 121 -499 1097
rect -275 121 -241 1097
rect -17 121 17 1097
rect 241 121 275 1097
rect 499 121 533 1097
rect 757 121 791 1097
rect 1015 121 1049 1097
rect 1273 121 1307 1097
rect 1531 121 1565 1097
rect 1789 121 1823 1097
rect 2047 121 2081 1097
rect 2305 121 2339 1097
rect 2563 121 2597 1097
rect 2821 121 2855 1097
rect 3079 121 3113 1097
rect 3337 121 3371 1097
rect 3595 121 3629 1097
rect -3629 -1097 -3595 -121
rect -3371 -1097 -3337 -121
rect -3113 -1097 -3079 -121
rect -2855 -1097 -2821 -121
rect -2597 -1097 -2563 -121
rect -2339 -1097 -2305 -121
rect -2081 -1097 -2047 -121
rect -1823 -1097 -1789 -121
rect -1565 -1097 -1531 -121
rect -1307 -1097 -1273 -121
rect -1049 -1097 -1015 -121
rect -791 -1097 -757 -121
rect -533 -1097 -499 -121
rect -275 -1097 -241 -121
rect -17 -1097 17 -121
rect 241 -1097 275 -121
rect 499 -1097 533 -121
rect 757 -1097 791 -121
rect 1015 -1097 1049 -121
rect 1273 -1097 1307 -121
rect 1531 -1097 1565 -121
rect 1789 -1097 1823 -121
rect 2047 -1097 2081 -121
rect 2305 -1097 2339 -121
rect 2563 -1097 2597 -121
rect 2821 -1097 2855 -121
rect 3079 -1097 3113 -121
rect 3337 -1097 3371 -121
rect 3595 -1097 3629 -121
<< mvpsubdiff >>
rect -3775 1319 3775 1331
rect -3775 1285 -3667 1319
rect 3667 1285 3775 1319
rect -3775 1273 3775 1285
rect -3775 1223 -3717 1273
rect -3775 -1223 -3763 1223
rect -3729 -1223 -3717 1223
rect 3717 1223 3775 1273
rect -3775 -1273 -3717 -1223
rect 3717 -1223 3729 1223
rect 3763 -1223 3775 1223
rect 3717 -1273 3775 -1223
rect -3775 -1285 3775 -1273
rect -3775 -1319 -3667 -1285
rect 3667 -1319 3775 -1285
rect -3775 -1331 3775 -1319
<< mvpsubdiffcont >>
rect -3667 1285 3667 1319
rect -3763 -1223 -3729 1223
rect 3729 -1223 3763 1223
rect -3667 -1319 3667 -1285
<< poly >>
rect -3583 1181 -3383 1197
rect -3583 1147 -3567 1181
rect -3399 1147 -3383 1181
rect -3583 1109 -3383 1147
rect -3325 1181 -3125 1197
rect -3325 1147 -3309 1181
rect -3141 1147 -3125 1181
rect -3325 1109 -3125 1147
rect -3067 1181 -2867 1197
rect -3067 1147 -3051 1181
rect -2883 1147 -2867 1181
rect -3067 1109 -2867 1147
rect -2809 1181 -2609 1197
rect -2809 1147 -2793 1181
rect -2625 1147 -2609 1181
rect -2809 1109 -2609 1147
rect -2551 1181 -2351 1197
rect -2551 1147 -2535 1181
rect -2367 1147 -2351 1181
rect -2551 1109 -2351 1147
rect -2293 1181 -2093 1197
rect -2293 1147 -2277 1181
rect -2109 1147 -2093 1181
rect -2293 1109 -2093 1147
rect -2035 1181 -1835 1197
rect -2035 1147 -2019 1181
rect -1851 1147 -1835 1181
rect -2035 1109 -1835 1147
rect -1777 1181 -1577 1197
rect -1777 1147 -1761 1181
rect -1593 1147 -1577 1181
rect -1777 1109 -1577 1147
rect -1519 1181 -1319 1197
rect -1519 1147 -1503 1181
rect -1335 1147 -1319 1181
rect -1519 1109 -1319 1147
rect -1261 1181 -1061 1197
rect -1261 1147 -1245 1181
rect -1077 1147 -1061 1181
rect -1261 1109 -1061 1147
rect -1003 1181 -803 1197
rect -1003 1147 -987 1181
rect -819 1147 -803 1181
rect -1003 1109 -803 1147
rect -745 1181 -545 1197
rect -745 1147 -729 1181
rect -561 1147 -545 1181
rect -745 1109 -545 1147
rect -487 1181 -287 1197
rect -487 1147 -471 1181
rect -303 1147 -287 1181
rect -487 1109 -287 1147
rect -229 1181 -29 1197
rect -229 1147 -213 1181
rect -45 1147 -29 1181
rect -229 1109 -29 1147
rect 29 1181 229 1197
rect 29 1147 45 1181
rect 213 1147 229 1181
rect 29 1109 229 1147
rect 287 1181 487 1197
rect 287 1147 303 1181
rect 471 1147 487 1181
rect 287 1109 487 1147
rect 545 1181 745 1197
rect 545 1147 561 1181
rect 729 1147 745 1181
rect 545 1109 745 1147
rect 803 1181 1003 1197
rect 803 1147 819 1181
rect 987 1147 1003 1181
rect 803 1109 1003 1147
rect 1061 1181 1261 1197
rect 1061 1147 1077 1181
rect 1245 1147 1261 1181
rect 1061 1109 1261 1147
rect 1319 1181 1519 1197
rect 1319 1147 1335 1181
rect 1503 1147 1519 1181
rect 1319 1109 1519 1147
rect 1577 1181 1777 1197
rect 1577 1147 1593 1181
rect 1761 1147 1777 1181
rect 1577 1109 1777 1147
rect 1835 1181 2035 1197
rect 1835 1147 1851 1181
rect 2019 1147 2035 1181
rect 1835 1109 2035 1147
rect 2093 1181 2293 1197
rect 2093 1147 2109 1181
rect 2277 1147 2293 1181
rect 2093 1109 2293 1147
rect 2351 1181 2551 1197
rect 2351 1147 2367 1181
rect 2535 1147 2551 1181
rect 2351 1109 2551 1147
rect 2609 1181 2809 1197
rect 2609 1147 2625 1181
rect 2793 1147 2809 1181
rect 2609 1109 2809 1147
rect 2867 1181 3067 1197
rect 2867 1147 2883 1181
rect 3051 1147 3067 1181
rect 2867 1109 3067 1147
rect 3125 1181 3325 1197
rect 3125 1147 3141 1181
rect 3309 1147 3325 1181
rect 3125 1109 3325 1147
rect 3383 1181 3583 1197
rect 3383 1147 3399 1181
rect 3567 1147 3583 1181
rect 3383 1109 3583 1147
rect -3583 71 -3383 109
rect -3583 37 -3567 71
rect -3399 37 -3383 71
rect -3583 21 -3383 37
rect -3325 71 -3125 109
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3325 21 -3125 37
rect -3067 71 -2867 109
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -3067 21 -2867 37
rect -2809 71 -2609 109
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2809 21 -2609 37
rect -2551 71 -2351 109
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2551 21 -2351 37
rect -2293 71 -2093 109
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2293 21 -2093 37
rect -2035 71 -1835 109
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 109
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 109
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 109
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 109
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 109
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 109
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 109
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect 2093 71 2293 109
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2093 21 2293 37
rect 2351 71 2551 109
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2351 21 2551 37
rect 2609 71 2809 109
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2609 21 2809 37
rect 2867 71 3067 109
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 2867 21 3067 37
rect 3125 71 3325 109
rect 3125 37 3141 71
rect 3309 37 3325 71
rect 3125 21 3325 37
rect 3383 71 3583 109
rect 3383 37 3399 71
rect 3567 37 3583 71
rect 3383 21 3583 37
rect -3583 -37 -3383 -21
rect -3583 -71 -3567 -37
rect -3399 -71 -3383 -37
rect -3583 -109 -3383 -71
rect -3325 -37 -3125 -21
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3325 -109 -3125 -71
rect -3067 -37 -2867 -21
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -3067 -109 -2867 -71
rect -2809 -37 -2609 -21
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2809 -109 -2609 -71
rect -2551 -37 -2351 -21
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2551 -109 -2351 -71
rect -2293 -37 -2093 -21
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2293 -109 -2093 -71
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -109 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -109 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -109 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -109 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -109 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -109 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -109 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -109 2035 -71
rect 2093 -37 2293 -21
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2093 -109 2293 -71
rect 2351 -37 2551 -21
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2351 -109 2551 -71
rect 2609 -37 2809 -21
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2609 -109 2809 -71
rect 2867 -37 3067 -21
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 2867 -109 3067 -71
rect 3125 -37 3325 -21
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect 3125 -109 3325 -71
rect 3383 -37 3583 -21
rect 3383 -71 3399 -37
rect 3567 -71 3583 -37
rect 3383 -109 3583 -71
rect -3583 -1147 -3383 -1109
rect -3583 -1181 -3567 -1147
rect -3399 -1181 -3383 -1147
rect -3583 -1197 -3383 -1181
rect -3325 -1147 -3125 -1109
rect -3325 -1181 -3309 -1147
rect -3141 -1181 -3125 -1147
rect -3325 -1197 -3125 -1181
rect -3067 -1147 -2867 -1109
rect -3067 -1181 -3051 -1147
rect -2883 -1181 -2867 -1147
rect -3067 -1197 -2867 -1181
rect -2809 -1147 -2609 -1109
rect -2809 -1181 -2793 -1147
rect -2625 -1181 -2609 -1147
rect -2809 -1197 -2609 -1181
rect -2551 -1147 -2351 -1109
rect -2551 -1181 -2535 -1147
rect -2367 -1181 -2351 -1147
rect -2551 -1197 -2351 -1181
rect -2293 -1147 -2093 -1109
rect -2293 -1181 -2277 -1147
rect -2109 -1181 -2093 -1147
rect -2293 -1197 -2093 -1181
rect -2035 -1147 -1835 -1109
rect -2035 -1181 -2019 -1147
rect -1851 -1181 -1835 -1147
rect -2035 -1197 -1835 -1181
rect -1777 -1147 -1577 -1109
rect -1777 -1181 -1761 -1147
rect -1593 -1181 -1577 -1147
rect -1777 -1197 -1577 -1181
rect -1519 -1147 -1319 -1109
rect -1519 -1181 -1503 -1147
rect -1335 -1181 -1319 -1147
rect -1519 -1197 -1319 -1181
rect -1261 -1147 -1061 -1109
rect -1261 -1181 -1245 -1147
rect -1077 -1181 -1061 -1147
rect -1261 -1197 -1061 -1181
rect -1003 -1147 -803 -1109
rect -1003 -1181 -987 -1147
rect -819 -1181 -803 -1147
rect -1003 -1197 -803 -1181
rect -745 -1147 -545 -1109
rect -745 -1181 -729 -1147
rect -561 -1181 -545 -1147
rect -745 -1197 -545 -1181
rect -487 -1147 -287 -1109
rect -487 -1181 -471 -1147
rect -303 -1181 -287 -1147
rect -487 -1197 -287 -1181
rect -229 -1147 -29 -1109
rect -229 -1181 -213 -1147
rect -45 -1181 -29 -1147
rect -229 -1197 -29 -1181
rect 29 -1147 229 -1109
rect 29 -1181 45 -1147
rect 213 -1181 229 -1147
rect 29 -1197 229 -1181
rect 287 -1147 487 -1109
rect 287 -1181 303 -1147
rect 471 -1181 487 -1147
rect 287 -1197 487 -1181
rect 545 -1147 745 -1109
rect 545 -1181 561 -1147
rect 729 -1181 745 -1147
rect 545 -1197 745 -1181
rect 803 -1147 1003 -1109
rect 803 -1181 819 -1147
rect 987 -1181 1003 -1147
rect 803 -1197 1003 -1181
rect 1061 -1147 1261 -1109
rect 1061 -1181 1077 -1147
rect 1245 -1181 1261 -1147
rect 1061 -1197 1261 -1181
rect 1319 -1147 1519 -1109
rect 1319 -1181 1335 -1147
rect 1503 -1181 1519 -1147
rect 1319 -1197 1519 -1181
rect 1577 -1147 1777 -1109
rect 1577 -1181 1593 -1147
rect 1761 -1181 1777 -1147
rect 1577 -1197 1777 -1181
rect 1835 -1147 2035 -1109
rect 1835 -1181 1851 -1147
rect 2019 -1181 2035 -1147
rect 1835 -1197 2035 -1181
rect 2093 -1147 2293 -1109
rect 2093 -1181 2109 -1147
rect 2277 -1181 2293 -1147
rect 2093 -1197 2293 -1181
rect 2351 -1147 2551 -1109
rect 2351 -1181 2367 -1147
rect 2535 -1181 2551 -1147
rect 2351 -1197 2551 -1181
rect 2609 -1147 2809 -1109
rect 2609 -1181 2625 -1147
rect 2793 -1181 2809 -1147
rect 2609 -1197 2809 -1181
rect 2867 -1147 3067 -1109
rect 2867 -1181 2883 -1147
rect 3051 -1181 3067 -1147
rect 2867 -1197 3067 -1181
rect 3125 -1147 3325 -1109
rect 3125 -1181 3141 -1147
rect 3309 -1181 3325 -1147
rect 3125 -1197 3325 -1181
rect 3383 -1147 3583 -1109
rect 3383 -1181 3399 -1147
rect 3567 -1181 3583 -1147
rect 3383 -1197 3583 -1181
<< polycont >>
rect -3567 1147 -3399 1181
rect -3309 1147 -3141 1181
rect -3051 1147 -2883 1181
rect -2793 1147 -2625 1181
rect -2535 1147 -2367 1181
rect -2277 1147 -2109 1181
rect -2019 1147 -1851 1181
rect -1761 1147 -1593 1181
rect -1503 1147 -1335 1181
rect -1245 1147 -1077 1181
rect -987 1147 -819 1181
rect -729 1147 -561 1181
rect -471 1147 -303 1181
rect -213 1147 -45 1181
rect 45 1147 213 1181
rect 303 1147 471 1181
rect 561 1147 729 1181
rect 819 1147 987 1181
rect 1077 1147 1245 1181
rect 1335 1147 1503 1181
rect 1593 1147 1761 1181
rect 1851 1147 2019 1181
rect 2109 1147 2277 1181
rect 2367 1147 2535 1181
rect 2625 1147 2793 1181
rect 2883 1147 3051 1181
rect 3141 1147 3309 1181
rect 3399 1147 3567 1181
rect -3567 37 -3399 71
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect 3399 37 3567 71
rect -3567 -71 -3399 -37
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect 3399 -71 3567 -37
rect -3567 -1181 -3399 -1147
rect -3309 -1181 -3141 -1147
rect -3051 -1181 -2883 -1147
rect -2793 -1181 -2625 -1147
rect -2535 -1181 -2367 -1147
rect -2277 -1181 -2109 -1147
rect -2019 -1181 -1851 -1147
rect -1761 -1181 -1593 -1147
rect -1503 -1181 -1335 -1147
rect -1245 -1181 -1077 -1147
rect -987 -1181 -819 -1147
rect -729 -1181 -561 -1147
rect -471 -1181 -303 -1147
rect -213 -1181 -45 -1147
rect 45 -1181 213 -1147
rect 303 -1181 471 -1147
rect 561 -1181 729 -1147
rect 819 -1181 987 -1147
rect 1077 -1181 1245 -1147
rect 1335 -1181 1503 -1147
rect 1593 -1181 1761 -1147
rect 1851 -1181 2019 -1147
rect 2109 -1181 2277 -1147
rect 2367 -1181 2535 -1147
rect 2625 -1181 2793 -1147
rect 2883 -1181 3051 -1147
rect 3141 -1181 3309 -1147
rect 3399 -1181 3567 -1147
<< locali >>
rect -3763 1285 -3667 1319
rect 3667 1285 3763 1319
rect -3763 1223 -3729 1285
rect 3729 1223 3763 1285
rect -3583 1147 -3567 1181
rect -3399 1147 -3383 1181
rect -3325 1147 -3309 1181
rect -3141 1147 -3125 1181
rect -3067 1147 -3051 1181
rect -2883 1147 -2867 1181
rect -2809 1147 -2793 1181
rect -2625 1147 -2609 1181
rect -2551 1147 -2535 1181
rect -2367 1147 -2351 1181
rect -2293 1147 -2277 1181
rect -2109 1147 -2093 1181
rect -2035 1147 -2019 1181
rect -1851 1147 -1835 1181
rect -1777 1147 -1761 1181
rect -1593 1147 -1577 1181
rect -1519 1147 -1503 1181
rect -1335 1147 -1319 1181
rect -1261 1147 -1245 1181
rect -1077 1147 -1061 1181
rect -1003 1147 -987 1181
rect -819 1147 -803 1181
rect -745 1147 -729 1181
rect -561 1147 -545 1181
rect -487 1147 -471 1181
rect -303 1147 -287 1181
rect -229 1147 -213 1181
rect -45 1147 -29 1181
rect 29 1147 45 1181
rect 213 1147 229 1181
rect 287 1147 303 1181
rect 471 1147 487 1181
rect 545 1147 561 1181
rect 729 1147 745 1181
rect 803 1147 819 1181
rect 987 1147 1003 1181
rect 1061 1147 1077 1181
rect 1245 1147 1261 1181
rect 1319 1147 1335 1181
rect 1503 1147 1519 1181
rect 1577 1147 1593 1181
rect 1761 1147 1777 1181
rect 1835 1147 1851 1181
rect 2019 1147 2035 1181
rect 2093 1147 2109 1181
rect 2277 1147 2293 1181
rect 2351 1147 2367 1181
rect 2535 1147 2551 1181
rect 2609 1147 2625 1181
rect 2793 1147 2809 1181
rect 2867 1147 2883 1181
rect 3051 1147 3067 1181
rect 3125 1147 3141 1181
rect 3309 1147 3325 1181
rect 3383 1147 3399 1181
rect 3567 1147 3583 1181
rect -3629 1097 -3595 1113
rect -3629 105 -3595 121
rect -3371 1097 -3337 1113
rect -3371 105 -3337 121
rect -3113 1097 -3079 1113
rect -3113 105 -3079 121
rect -2855 1097 -2821 1113
rect -2855 105 -2821 121
rect -2597 1097 -2563 1113
rect -2597 105 -2563 121
rect -2339 1097 -2305 1113
rect -2339 105 -2305 121
rect -2081 1097 -2047 1113
rect -2081 105 -2047 121
rect -1823 1097 -1789 1113
rect -1823 105 -1789 121
rect -1565 1097 -1531 1113
rect -1565 105 -1531 121
rect -1307 1097 -1273 1113
rect -1307 105 -1273 121
rect -1049 1097 -1015 1113
rect -1049 105 -1015 121
rect -791 1097 -757 1113
rect -791 105 -757 121
rect -533 1097 -499 1113
rect -533 105 -499 121
rect -275 1097 -241 1113
rect -275 105 -241 121
rect -17 1097 17 1113
rect -17 105 17 121
rect 241 1097 275 1113
rect 241 105 275 121
rect 499 1097 533 1113
rect 499 105 533 121
rect 757 1097 791 1113
rect 757 105 791 121
rect 1015 1097 1049 1113
rect 1015 105 1049 121
rect 1273 1097 1307 1113
rect 1273 105 1307 121
rect 1531 1097 1565 1113
rect 1531 105 1565 121
rect 1789 1097 1823 1113
rect 1789 105 1823 121
rect 2047 1097 2081 1113
rect 2047 105 2081 121
rect 2305 1097 2339 1113
rect 2305 105 2339 121
rect 2563 1097 2597 1113
rect 2563 105 2597 121
rect 2821 1097 2855 1113
rect 2821 105 2855 121
rect 3079 1097 3113 1113
rect 3079 105 3113 121
rect 3337 1097 3371 1113
rect 3337 105 3371 121
rect 3595 1097 3629 1113
rect 3595 105 3629 121
rect -3583 37 -3567 71
rect -3399 37 -3383 71
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 3125 37 3141 71
rect 3309 37 3325 71
rect 3383 37 3399 71
rect 3567 37 3583 71
rect -3583 -71 -3567 -37
rect -3399 -71 -3383 -37
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect 3383 -71 3399 -37
rect 3567 -71 3583 -37
rect -3629 -121 -3595 -105
rect -3629 -1113 -3595 -1097
rect -3371 -121 -3337 -105
rect -3371 -1113 -3337 -1097
rect -3113 -121 -3079 -105
rect -3113 -1113 -3079 -1097
rect -2855 -121 -2821 -105
rect -2855 -1113 -2821 -1097
rect -2597 -121 -2563 -105
rect -2597 -1113 -2563 -1097
rect -2339 -121 -2305 -105
rect -2339 -1113 -2305 -1097
rect -2081 -121 -2047 -105
rect -2081 -1113 -2047 -1097
rect -1823 -121 -1789 -105
rect -1823 -1113 -1789 -1097
rect -1565 -121 -1531 -105
rect -1565 -1113 -1531 -1097
rect -1307 -121 -1273 -105
rect -1307 -1113 -1273 -1097
rect -1049 -121 -1015 -105
rect -1049 -1113 -1015 -1097
rect -791 -121 -757 -105
rect -791 -1113 -757 -1097
rect -533 -121 -499 -105
rect -533 -1113 -499 -1097
rect -275 -121 -241 -105
rect -275 -1113 -241 -1097
rect -17 -121 17 -105
rect -17 -1113 17 -1097
rect 241 -121 275 -105
rect 241 -1113 275 -1097
rect 499 -121 533 -105
rect 499 -1113 533 -1097
rect 757 -121 791 -105
rect 757 -1113 791 -1097
rect 1015 -121 1049 -105
rect 1015 -1113 1049 -1097
rect 1273 -121 1307 -105
rect 1273 -1113 1307 -1097
rect 1531 -121 1565 -105
rect 1531 -1113 1565 -1097
rect 1789 -121 1823 -105
rect 1789 -1113 1823 -1097
rect 2047 -121 2081 -105
rect 2047 -1113 2081 -1097
rect 2305 -121 2339 -105
rect 2305 -1113 2339 -1097
rect 2563 -121 2597 -105
rect 2563 -1113 2597 -1097
rect 2821 -121 2855 -105
rect 2821 -1113 2855 -1097
rect 3079 -121 3113 -105
rect 3079 -1113 3113 -1097
rect 3337 -121 3371 -105
rect 3337 -1113 3371 -1097
rect 3595 -121 3629 -105
rect 3595 -1113 3629 -1097
rect -3583 -1181 -3567 -1147
rect -3399 -1181 -3383 -1147
rect -3325 -1181 -3309 -1147
rect -3141 -1181 -3125 -1147
rect -3067 -1181 -3051 -1147
rect -2883 -1181 -2867 -1147
rect -2809 -1181 -2793 -1147
rect -2625 -1181 -2609 -1147
rect -2551 -1181 -2535 -1147
rect -2367 -1181 -2351 -1147
rect -2293 -1181 -2277 -1147
rect -2109 -1181 -2093 -1147
rect -2035 -1181 -2019 -1147
rect -1851 -1181 -1835 -1147
rect -1777 -1181 -1761 -1147
rect -1593 -1181 -1577 -1147
rect -1519 -1181 -1503 -1147
rect -1335 -1181 -1319 -1147
rect -1261 -1181 -1245 -1147
rect -1077 -1181 -1061 -1147
rect -1003 -1181 -987 -1147
rect -819 -1181 -803 -1147
rect -745 -1181 -729 -1147
rect -561 -1181 -545 -1147
rect -487 -1181 -471 -1147
rect -303 -1181 -287 -1147
rect -229 -1181 -213 -1147
rect -45 -1181 -29 -1147
rect 29 -1181 45 -1147
rect 213 -1181 229 -1147
rect 287 -1181 303 -1147
rect 471 -1181 487 -1147
rect 545 -1181 561 -1147
rect 729 -1181 745 -1147
rect 803 -1181 819 -1147
rect 987 -1181 1003 -1147
rect 1061 -1181 1077 -1147
rect 1245 -1181 1261 -1147
rect 1319 -1181 1335 -1147
rect 1503 -1181 1519 -1147
rect 1577 -1181 1593 -1147
rect 1761 -1181 1777 -1147
rect 1835 -1181 1851 -1147
rect 2019 -1181 2035 -1147
rect 2093 -1181 2109 -1147
rect 2277 -1181 2293 -1147
rect 2351 -1181 2367 -1147
rect 2535 -1181 2551 -1147
rect 2609 -1181 2625 -1147
rect 2793 -1181 2809 -1147
rect 2867 -1181 2883 -1147
rect 3051 -1181 3067 -1147
rect 3125 -1181 3141 -1147
rect 3309 -1181 3325 -1147
rect 3383 -1181 3399 -1147
rect 3567 -1181 3583 -1147
rect -3763 -1285 -3729 -1223
rect 3729 -1285 3763 -1223
rect -3763 -1319 -3667 -1285
rect 3667 -1319 3763 -1285
<< viali >>
rect -3567 1147 -3399 1181
rect -3309 1147 -3141 1181
rect -3051 1147 -2883 1181
rect -2793 1147 -2625 1181
rect -2535 1147 -2367 1181
rect -2277 1147 -2109 1181
rect -2019 1147 -1851 1181
rect -1761 1147 -1593 1181
rect -1503 1147 -1335 1181
rect -1245 1147 -1077 1181
rect -987 1147 -819 1181
rect -729 1147 -561 1181
rect -471 1147 -303 1181
rect -213 1147 -45 1181
rect 45 1147 213 1181
rect 303 1147 471 1181
rect 561 1147 729 1181
rect 819 1147 987 1181
rect 1077 1147 1245 1181
rect 1335 1147 1503 1181
rect 1593 1147 1761 1181
rect 1851 1147 2019 1181
rect 2109 1147 2277 1181
rect 2367 1147 2535 1181
rect 2625 1147 2793 1181
rect 2883 1147 3051 1181
rect 3141 1147 3309 1181
rect 3399 1147 3567 1181
rect -3629 121 -3595 1097
rect -3371 121 -3337 1097
rect -3113 121 -3079 1097
rect -2855 121 -2821 1097
rect -2597 121 -2563 1097
rect -2339 121 -2305 1097
rect -2081 121 -2047 1097
rect -1823 121 -1789 1097
rect -1565 121 -1531 1097
rect -1307 121 -1273 1097
rect -1049 121 -1015 1097
rect -791 121 -757 1097
rect -533 121 -499 1097
rect -275 121 -241 1097
rect -17 121 17 1097
rect 241 121 275 1097
rect 499 121 533 1097
rect 757 121 791 1097
rect 1015 121 1049 1097
rect 1273 121 1307 1097
rect 1531 121 1565 1097
rect 1789 121 1823 1097
rect 2047 121 2081 1097
rect 2305 121 2339 1097
rect 2563 121 2597 1097
rect 2821 121 2855 1097
rect 3079 121 3113 1097
rect 3337 121 3371 1097
rect 3595 121 3629 1097
rect -3567 37 -3399 71
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect 3399 37 3567 71
rect -3567 -71 -3399 -37
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect 3399 -71 3567 -37
rect -3629 -1097 -3595 -121
rect -3371 -1097 -3337 -121
rect -3113 -1097 -3079 -121
rect -2855 -1097 -2821 -121
rect -2597 -1097 -2563 -121
rect -2339 -1097 -2305 -121
rect -2081 -1097 -2047 -121
rect -1823 -1097 -1789 -121
rect -1565 -1097 -1531 -121
rect -1307 -1097 -1273 -121
rect -1049 -1097 -1015 -121
rect -791 -1097 -757 -121
rect -533 -1097 -499 -121
rect -275 -1097 -241 -121
rect -17 -1097 17 -121
rect 241 -1097 275 -121
rect 499 -1097 533 -121
rect 757 -1097 791 -121
rect 1015 -1097 1049 -121
rect 1273 -1097 1307 -121
rect 1531 -1097 1565 -121
rect 1789 -1097 1823 -121
rect 2047 -1097 2081 -121
rect 2305 -1097 2339 -121
rect 2563 -1097 2597 -121
rect 2821 -1097 2855 -121
rect 3079 -1097 3113 -121
rect 3337 -1097 3371 -121
rect 3595 -1097 3629 -121
rect -3567 -1181 -3399 -1147
rect -3309 -1181 -3141 -1147
rect -3051 -1181 -2883 -1147
rect -2793 -1181 -2625 -1147
rect -2535 -1181 -2367 -1147
rect -2277 -1181 -2109 -1147
rect -2019 -1181 -1851 -1147
rect -1761 -1181 -1593 -1147
rect -1503 -1181 -1335 -1147
rect -1245 -1181 -1077 -1147
rect -987 -1181 -819 -1147
rect -729 -1181 -561 -1147
rect -471 -1181 -303 -1147
rect -213 -1181 -45 -1147
rect 45 -1181 213 -1147
rect 303 -1181 471 -1147
rect 561 -1181 729 -1147
rect 819 -1181 987 -1147
rect 1077 -1181 1245 -1147
rect 1335 -1181 1503 -1147
rect 1593 -1181 1761 -1147
rect 1851 -1181 2019 -1147
rect 2109 -1181 2277 -1147
rect 2367 -1181 2535 -1147
rect 2625 -1181 2793 -1147
rect 2883 -1181 3051 -1147
rect 3141 -1181 3309 -1147
rect 3399 -1181 3567 -1147
<< metal1 >>
rect -3579 1181 -3387 1187
rect -3579 1147 -3567 1181
rect -3399 1147 -3387 1181
rect -3579 1141 -3387 1147
rect -3321 1181 -3129 1187
rect -3321 1147 -3309 1181
rect -3141 1147 -3129 1181
rect -3321 1141 -3129 1147
rect -3063 1181 -2871 1187
rect -3063 1147 -3051 1181
rect -2883 1147 -2871 1181
rect -3063 1141 -2871 1147
rect -2805 1181 -2613 1187
rect -2805 1147 -2793 1181
rect -2625 1147 -2613 1181
rect -2805 1141 -2613 1147
rect -2547 1181 -2355 1187
rect -2547 1147 -2535 1181
rect -2367 1147 -2355 1181
rect -2547 1141 -2355 1147
rect -2289 1181 -2097 1187
rect -2289 1147 -2277 1181
rect -2109 1147 -2097 1181
rect -2289 1141 -2097 1147
rect -2031 1181 -1839 1187
rect -2031 1147 -2019 1181
rect -1851 1147 -1839 1181
rect -2031 1141 -1839 1147
rect -1773 1181 -1581 1187
rect -1773 1147 -1761 1181
rect -1593 1147 -1581 1181
rect -1773 1141 -1581 1147
rect -1515 1181 -1323 1187
rect -1515 1147 -1503 1181
rect -1335 1147 -1323 1181
rect -1515 1141 -1323 1147
rect -1257 1181 -1065 1187
rect -1257 1147 -1245 1181
rect -1077 1147 -1065 1181
rect -1257 1141 -1065 1147
rect -999 1181 -807 1187
rect -999 1147 -987 1181
rect -819 1147 -807 1181
rect -999 1141 -807 1147
rect -741 1181 -549 1187
rect -741 1147 -729 1181
rect -561 1147 -549 1181
rect -741 1141 -549 1147
rect -483 1181 -291 1187
rect -483 1147 -471 1181
rect -303 1147 -291 1181
rect -483 1141 -291 1147
rect -225 1181 -33 1187
rect -225 1147 -213 1181
rect -45 1147 -33 1181
rect -225 1141 -33 1147
rect 33 1181 225 1187
rect 33 1147 45 1181
rect 213 1147 225 1181
rect 33 1141 225 1147
rect 291 1181 483 1187
rect 291 1147 303 1181
rect 471 1147 483 1181
rect 291 1141 483 1147
rect 549 1181 741 1187
rect 549 1147 561 1181
rect 729 1147 741 1181
rect 549 1141 741 1147
rect 807 1181 999 1187
rect 807 1147 819 1181
rect 987 1147 999 1181
rect 807 1141 999 1147
rect 1065 1181 1257 1187
rect 1065 1147 1077 1181
rect 1245 1147 1257 1181
rect 1065 1141 1257 1147
rect 1323 1181 1515 1187
rect 1323 1147 1335 1181
rect 1503 1147 1515 1181
rect 1323 1141 1515 1147
rect 1581 1181 1773 1187
rect 1581 1147 1593 1181
rect 1761 1147 1773 1181
rect 1581 1141 1773 1147
rect 1839 1181 2031 1187
rect 1839 1147 1851 1181
rect 2019 1147 2031 1181
rect 1839 1141 2031 1147
rect 2097 1181 2289 1187
rect 2097 1147 2109 1181
rect 2277 1147 2289 1181
rect 2097 1141 2289 1147
rect 2355 1181 2547 1187
rect 2355 1147 2367 1181
rect 2535 1147 2547 1181
rect 2355 1141 2547 1147
rect 2613 1181 2805 1187
rect 2613 1147 2625 1181
rect 2793 1147 2805 1181
rect 2613 1141 2805 1147
rect 2871 1181 3063 1187
rect 2871 1147 2883 1181
rect 3051 1147 3063 1181
rect 2871 1141 3063 1147
rect 3129 1181 3321 1187
rect 3129 1147 3141 1181
rect 3309 1147 3321 1181
rect 3129 1141 3321 1147
rect 3387 1181 3579 1187
rect 3387 1147 3399 1181
rect 3567 1147 3579 1181
rect 3387 1141 3579 1147
rect -3635 1097 -3589 1109
rect -3635 121 -3629 1097
rect -3595 121 -3589 1097
rect -3635 109 -3589 121
rect -3377 1097 -3331 1109
rect -3377 121 -3371 1097
rect -3337 121 -3331 1097
rect -3377 109 -3331 121
rect -3119 1097 -3073 1109
rect -3119 121 -3113 1097
rect -3079 121 -3073 1097
rect -3119 109 -3073 121
rect -2861 1097 -2815 1109
rect -2861 121 -2855 1097
rect -2821 121 -2815 1097
rect -2861 109 -2815 121
rect -2603 1097 -2557 1109
rect -2603 121 -2597 1097
rect -2563 121 -2557 1097
rect -2603 109 -2557 121
rect -2345 1097 -2299 1109
rect -2345 121 -2339 1097
rect -2305 121 -2299 1097
rect -2345 109 -2299 121
rect -2087 1097 -2041 1109
rect -2087 121 -2081 1097
rect -2047 121 -2041 1097
rect -2087 109 -2041 121
rect -1829 1097 -1783 1109
rect -1829 121 -1823 1097
rect -1789 121 -1783 1097
rect -1829 109 -1783 121
rect -1571 1097 -1525 1109
rect -1571 121 -1565 1097
rect -1531 121 -1525 1097
rect -1571 109 -1525 121
rect -1313 1097 -1267 1109
rect -1313 121 -1307 1097
rect -1273 121 -1267 1097
rect -1313 109 -1267 121
rect -1055 1097 -1009 1109
rect -1055 121 -1049 1097
rect -1015 121 -1009 1097
rect -1055 109 -1009 121
rect -797 1097 -751 1109
rect -797 121 -791 1097
rect -757 121 -751 1097
rect -797 109 -751 121
rect -539 1097 -493 1109
rect -539 121 -533 1097
rect -499 121 -493 1097
rect -539 109 -493 121
rect -281 1097 -235 1109
rect -281 121 -275 1097
rect -241 121 -235 1097
rect -281 109 -235 121
rect -23 1097 23 1109
rect -23 121 -17 1097
rect 17 121 23 1097
rect -23 109 23 121
rect 235 1097 281 1109
rect 235 121 241 1097
rect 275 121 281 1097
rect 235 109 281 121
rect 493 1097 539 1109
rect 493 121 499 1097
rect 533 121 539 1097
rect 493 109 539 121
rect 751 1097 797 1109
rect 751 121 757 1097
rect 791 121 797 1097
rect 751 109 797 121
rect 1009 1097 1055 1109
rect 1009 121 1015 1097
rect 1049 121 1055 1097
rect 1009 109 1055 121
rect 1267 1097 1313 1109
rect 1267 121 1273 1097
rect 1307 121 1313 1097
rect 1267 109 1313 121
rect 1525 1097 1571 1109
rect 1525 121 1531 1097
rect 1565 121 1571 1097
rect 1525 109 1571 121
rect 1783 1097 1829 1109
rect 1783 121 1789 1097
rect 1823 121 1829 1097
rect 1783 109 1829 121
rect 2041 1097 2087 1109
rect 2041 121 2047 1097
rect 2081 121 2087 1097
rect 2041 109 2087 121
rect 2299 1097 2345 1109
rect 2299 121 2305 1097
rect 2339 121 2345 1097
rect 2299 109 2345 121
rect 2557 1097 2603 1109
rect 2557 121 2563 1097
rect 2597 121 2603 1097
rect 2557 109 2603 121
rect 2815 1097 2861 1109
rect 2815 121 2821 1097
rect 2855 121 2861 1097
rect 2815 109 2861 121
rect 3073 1097 3119 1109
rect 3073 121 3079 1097
rect 3113 121 3119 1097
rect 3073 109 3119 121
rect 3331 1097 3377 1109
rect 3331 121 3337 1097
rect 3371 121 3377 1097
rect 3331 109 3377 121
rect 3589 1097 3635 1109
rect 3589 121 3595 1097
rect 3629 121 3635 1097
rect 3589 109 3635 121
rect -3579 71 -3387 77
rect -3579 37 -3567 71
rect -3399 37 -3387 71
rect -3579 31 -3387 37
rect -3321 71 -3129 77
rect -3321 37 -3309 71
rect -3141 37 -3129 71
rect -3321 31 -3129 37
rect -3063 71 -2871 77
rect -3063 37 -3051 71
rect -2883 37 -2871 71
rect -3063 31 -2871 37
rect -2805 71 -2613 77
rect -2805 37 -2793 71
rect -2625 37 -2613 71
rect -2805 31 -2613 37
rect -2547 71 -2355 77
rect -2547 37 -2535 71
rect -2367 37 -2355 71
rect -2547 31 -2355 37
rect -2289 71 -2097 77
rect -2289 37 -2277 71
rect -2109 37 -2097 71
rect -2289 31 -2097 37
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect 2097 71 2289 77
rect 2097 37 2109 71
rect 2277 37 2289 71
rect 2097 31 2289 37
rect 2355 71 2547 77
rect 2355 37 2367 71
rect 2535 37 2547 71
rect 2355 31 2547 37
rect 2613 71 2805 77
rect 2613 37 2625 71
rect 2793 37 2805 71
rect 2613 31 2805 37
rect 2871 71 3063 77
rect 2871 37 2883 71
rect 3051 37 3063 71
rect 2871 31 3063 37
rect 3129 71 3321 77
rect 3129 37 3141 71
rect 3309 37 3321 71
rect 3129 31 3321 37
rect 3387 71 3579 77
rect 3387 37 3399 71
rect 3567 37 3579 71
rect 3387 31 3579 37
rect -3579 -37 -3387 -31
rect -3579 -71 -3567 -37
rect -3399 -71 -3387 -37
rect -3579 -77 -3387 -71
rect -3321 -37 -3129 -31
rect -3321 -71 -3309 -37
rect -3141 -71 -3129 -37
rect -3321 -77 -3129 -71
rect -3063 -37 -2871 -31
rect -3063 -71 -3051 -37
rect -2883 -71 -2871 -37
rect -3063 -77 -2871 -71
rect -2805 -37 -2613 -31
rect -2805 -71 -2793 -37
rect -2625 -71 -2613 -37
rect -2805 -77 -2613 -71
rect -2547 -37 -2355 -31
rect -2547 -71 -2535 -37
rect -2367 -71 -2355 -37
rect -2547 -77 -2355 -71
rect -2289 -37 -2097 -31
rect -2289 -71 -2277 -37
rect -2109 -71 -2097 -37
rect -2289 -77 -2097 -71
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect 2097 -37 2289 -31
rect 2097 -71 2109 -37
rect 2277 -71 2289 -37
rect 2097 -77 2289 -71
rect 2355 -37 2547 -31
rect 2355 -71 2367 -37
rect 2535 -71 2547 -37
rect 2355 -77 2547 -71
rect 2613 -37 2805 -31
rect 2613 -71 2625 -37
rect 2793 -71 2805 -37
rect 2613 -77 2805 -71
rect 2871 -37 3063 -31
rect 2871 -71 2883 -37
rect 3051 -71 3063 -37
rect 2871 -77 3063 -71
rect 3129 -37 3321 -31
rect 3129 -71 3141 -37
rect 3309 -71 3321 -37
rect 3129 -77 3321 -71
rect 3387 -37 3579 -31
rect 3387 -71 3399 -37
rect 3567 -71 3579 -37
rect 3387 -77 3579 -71
rect -3635 -121 -3589 -109
rect -3635 -1097 -3629 -121
rect -3595 -1097 -3589 -121
rect -3635 -1109 -3589 -1097
rect -3377 -121 -3331 -109
rect -3377 -1097 -3371 -121
rect -3337 -1097 -3331 -121
rect -3377 -1109 -3331 -1097
rect -3119 -121 -3073 -109
rect -3119 -1097 -3113 -121
rect -3079 -1097 -3073 -121
rect -3119 -1109 -3073 -1097
rect -2861 -121 -2815 -109
rect -2861 -1097 -2855 -121
rect -2821 -1097 -2815 -121
rect -2861 -1109 -2815 -1097
rect -2603 -121 -2557 -109
rect -2603 -1097 -2597 -121
rect -2563 -1097 -2557 -121
rect -2603 -1109 -2557 -1097
rect -2345 -121 -2299 -109
rect -2345 -1097 -2339 -121
rect -2305 -1097 -2299 -121
rect -2345 -1109 -2299 -1097
rect -2087 -121 -2041 -109
rect -2087 -1097 -2081 -121
rect -2047 -1097 -2041 -121
rect -2087 -1109 -2041 -1097
rect -1829 -121 -1783 -109
rect -1829 -1097 -1823 -121
rect -1789 -1097 -1783 -121
rect -1829 -1109 -1783 -1097
rect -1571 -121 -1525 -109
rect -1571 -1097 -1565 -121
rect -1531 -1097 -1525 -121
rect -1571 -1109 -1525 -1097
rect -1313 -121 -1267 -109
rect -1313 -1097 -1307 -121
rect -1273 -1097 -1267 -121
rect -1313 -1109 -1267 -1097
rect -1055 -121 -1009 -109
rect -1055 -1097 -1049 -121
rect -1015 -1097 -1009 -121
rect -1055 -1109 -1009 -1097
rect -797 -121 -751 -109
rect -797 -1097 -791 -121
rect -757 -1097 -751 -121
rect -797 -1109 -751 -1097
rect -539 -121 -493 -109
rect -539 -1097 -533 -121
rect -499 -1097 -493 -121
rect -539 -1109 -493 -1097
rect -281 -121 -235 -109
rect -281 -1097 -275 -121
rect -241 -1097 -235 -121
rect -281 -1109 -235 -1097
rect -23 -121 23 -109
rect -23 -1097 -17 -121
rect 17 -1097 23 -121
rect -23 -1109 23 -1097
rect 235 -121 281 -109
rect 235 -1097 241 -121
rect 275 -1097 281 -121
rect 235 -1109 281 -1097
rect 493 -121 539 -109
rect 493 -1097 499 -121
rect 533 -1097 539 -121
rect 493 -1109 539 -1097
rect 751 -121 797 -109
rect 751 -1097 757 -121
rect 791 -1097 797 -121
rect 751 -1109 797 -1097
rect 1009 -121 1055 -109
rect 1009 -1097 1015 -121
rect 1049 -1097 1055 -121
rect 1009 -1109 1055 -1097
rect 1267 -121 1313 -109
rect 1267 -1097 1273 -121
rect 1307 -1097 1313 -121
rect 1267 -1109 1313 -1097
rect 1525 -121 1571 -109
rect 1525 -1097 1531 -121
rect 1565 -1097 1571 -121
rect 1525 -1109 1571 -1097
rect 1783 -121 1829 -109
rect 1783 -1097 1789 -121
rect 1823 -1097 1829 -121
rect 1783 -1109 1829 -1097
rect 2041 -121 2087 -109
rect 2041 -1097 2047 -121
rect 2081 -1097 2087 -121
rect 2041 -1109 2087 -1097
rect 2299 -121 2345 -109
rect 2299 -1097 2305 -121
rect 2339 -1097 2345 -121
rect 2299 -1109 2345 -1097
rect 2557 -121 2603 -109
rect 2557 -1097 2563 -121
rect 2597 -1097 2603 -121
rect 2557 -1109 2603 -1097
rect 2815 -121 2861 -109
rect 2815 -1097 2821 -121
rect 2855 -1097 2861 -121
rect 2815 -1109 2861 -1097
rect 3073 -121 3119 -109
rect 3073 -1097 3079 -121
rect 3113 -1097 3119 -121
rect 3073 -1109 3119 -1097
rect 3331 -121 3377 -109
rect 3331 -1097 3337 -121
rect 3371 -1097 3377 -121
rect 3331 -1109 3377 -1097
rect 3589 -121 3635 -109
rect 3589 -1097 3595 -121
rect 3629 -1097 3635 -121
rect 3589 -1109 3635 -1097
rect -3579 -1147 -3387 -1141
rect -3579 -1181 -3567 -1147
rect -3399 -1181 -3387 -1147
rect -3579 -1187 -3387 -1181
rect -3321 -1147 -3129 -1141
rect -3321 -1181 -3309 -1147
rect -3141 -1181 -3129 -1147
rect -3321 -1187 -3129 -1181
rect -3063 -1147 -2871 -1141
rect -3063 -1181 -3051 -1147
rect -2883 -1181 -2871 -1147
rect -3063 -1187 -2871 -1181
rect -2805 -1147 -2613 -1141
rect -2805 -1181 -2793 -1147
rect -2625 -1181 -2613 -1147
rect -2805 -1187 -2613 -1181
rect -2547 -1147 -2355 -1141
rect -2547 -1181 -2535 -1147
rect -2367 -1181 -2355 -1147
rect -2547 -1187 -2355 -1181
rect -2289 -1147 -2097 -1141
rect -2289 -1181 -2277 -1147
rect -2109 -1181 -2097 -1147
rect -2289 -1187 -2097 -1181
rect -2031 -1147 -1839 -1141
rect -2031 -1181 -2019 -1147
rect -1851 -1181 -1839 -1147
rect -2031 -1187 -1839 -1181
rect -1773 -1147 -1581 -1141
rect -1773 -1181 -1761 -1147
rect -1593 -1181 -1581 -1147
rect -1773 -1187 -1581 -1181
rect -1515 -1147 -1323 -1141
rect -1515 -1181 -1503 -1147
rect -1335 -1181 -1323 -1147
rect -1515 -1187 -1323 -1181
rect -1257 -1147 -1065 -1141
rect -1257 -1181 -1245 -1147
rect -1077 -1181 -1065 -1147
rect -1257 -1187 -1065 -1181
rect -999 -1147 -807 -1141
rect -999 -1181 -987 -1147
rect -819 -1181 -807 -1147
rect -999 -1187 -807 -1181
rect -741 -1147 -549 -1141
rect -741 -1181 -729 -1147
rect -561 -1181 -549 -1147
rect -741 -1187 -549 -1181
rect -483 -1147 -291 -1141
rect -483 -1181 -471 -1147
rect -303 -1181 -291 -1147
rect -483 -1187 -291 -1181
rect -225 -1147 -33 -1141
rect -225 -1181 -213 -1147
rect -45 -1181 -33 -1147
rect -225 -1187 -33 -1181
rect 33 -1147 225 -1141
rect 33 -1181 45 -1147
rect 213 -1181 225 -1147
rect 33 -1187 225 -1181
rect 291 -1147 483 -1141
rect 291 -1181 303 -1147
rect 471 -1181 483 -1147
rect 291 -1187 483 -1181
rect 549 -1147 741 -1141
rect 549 -1181 561 -1147
rect 729 -1181 741 -1147
rect 549 -1187 741 -1181
rect 807 -1147 999 -1141
rect 807 -1181 819 -1147
rect 987 -1181 999 -1147
rect 807 -1187 999 -1181
rect 1065 -1147 1257 -1141
rect 1065 -1181 1077 -1147
rect 1245 -1181 1257 -1147
rect 1065 -1187 1257 -1181
rect 1323 -1147 1515 -1141
rect 1323 -1181 1335 -1147
rect 1503 -1181 1515 -1147
rect 1323 -1187 1515 -1181
rect 1581 -1147 1773 -1141
rect 1581 -1181 1593 -1147
rect 1761 -1181 1773 -1147
rect 1581 -1187 1773 -1181
rect 1839 -1147 2031 -1141
rect 1839 -1181 1851 -1147
rect 2019 -1181 2031 -1147
rect 1839 -1187 2031 -1181
rect 2097 -1147 2289 -1141
rect 2097 -1181 2109 -1147
rect 2277 -1181 2289 -1147
rect 2097 -1187 2289 -1181
rect 2355 -1147 2547 -1141
rect 2355 -1181 2367 -1147
rect 2535 -1181 2547 -1147
rect 2355 -1187 2547 -1181
rect 2613 -1147 2805 -1141
rect 2613 -1181 2625 -1147
rect 2793 -1181 2805 -1147
rect 2613 -1187 2805 -1181
rect 2871 -1147 3063 -1141
rect 2871 -1181 2883 -1147
rect 3051 -1181 3063 -1147
rect 2871 -1187 3063 -1181
rect 3129 -1147 3321 -1141
rect 3129 -1181 3141 -1147
rect 3309 -1181 3321 -1147
rect 3129 -1187 3321 -1181
rect 3387 -1147 3579 -1141
rect 3387 -1181 3399 -1147
rect 3567 -1181 3579 -1147
rect 3387 -1187 3579 -1181
<< properties >>
string FIXED_BBOX -3746 -1302 3746 1302
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 2 nf 28 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1757785414
<< nwell >>
rect -2035 -1415 2035 1415
<< mvpmos >>
rect -1777 118 -1577 1118
rect -1519 118 -1319 1118
rect -1261 118 -1061 1118
rect -1003 118 -803 1118
rect -745 118 -545 1118
rect -487 118 -287 1118
rect -229 118 -29 1118
rect 29 118 229 1118
rect 287 118 487 1118
rect 545 118 745 1118
rect 803 118 1003 1118
rect 1061 118 1261 1118
rect 1319 118 1519 1118
rect 1577 118 1777 1118
rect -1777 -1118 -1577 -118
rect -1519 -1118 -1319 -118
rect -1261 -1118 -1061 -118
rect -1003 -1118 -803 -118
rect -745 -1118 -545 -118
rect -487 -1118 -287 -118
rect -229 -1118 -29 -118
rect 29 -1118 229 -118
rect 287 -1118 487 -118
rect 545 -1118 745 -118
rect 803 -1118 1003 -118
rect 1061 -1118 1261 -118
rect 1319 -1118 1519 -118
rect 1577 -1118 1777 -118
<< mvpdiff >>
rect -1835 1106 -1777 1118
rect -1835 130 -1823 1106
rect -1789 130 -1777 1106
rect -1835 118 -1777 130
rect -1577 1106 -1519 1118
rect -1577 130 -1565 1106
rect -1531 130 -1519 1106
rect -1577 118 -1519 130
rect -1319 1106 -1261 1118
rect -1319 130 -1307 1106
rect -1273 130 -1261 1106
rect -1319 118 -1261 130
rect -1061 1106 -1003 1118
rect -1061 130 -1049 1106
rect -1015 130 -1003 1106
rect -1061 118 -1003 130
rect -803 1106 -745 1118
rect -803 130 -791 1106
rect -757 130 -745 1106
rect -803 118 -745 130
rect -545 1106 -487 1118
rect -545 130 -533 1106
rect -499 130 -487 1106
rect -545 118 -487 130
rect -287 1106 -229 1118
rect -287 130 -275 1106
rect -241 130 -229 1106
rect -287 118 -229 130
rect -29 1106 29 1118
rect -29 130 -17 1106
rect 17 130 29 1106
rect -29 118 29 130
rect 229 1106 287 1118
rect 229 130 241 1106
rect 275 130 287 1106
rect 229 118 287 130
rect 487 1106 545 1118
rect 487 130 499 1106
rect 533 130 545 1106
rect 487 118 545 130
rect 745 1106 803 1118
rect 745 130 757 1106
rect 791 130 803 1106
rect 745 118 803 130
rect 1003 1106 1061 1118
rect 1003 130 1015 1106
rect 1049 130 1061 1106
rect 1003 118 1061 130
rect 1261 1106 1319 1118
rect 1261 130 1273 1106
rect 1307 130 1319 1106
rect 1261 118 1319 130
rect 1519 1106 1577 1118
rect 1519 130 1531 1106
rect 1565 130 1577 1106
rect 1519 118 1577 130
rect 1777 1106 1835 1118
rect 1777 130 1789 1106
rect 1823 130 1835 1106
rect 1777 118 1835 130
rect -1835 -130 -1777 -118
rect -1835 -1106 -1823 -130
rect -1789 -1106 -1777 -130
rect -1835 -1118 -1777 -1106
rect -1577 -130 -1519 -118
rect -1577 -1106 -1565 -130
rect -1531 -1106 -1519 -130
rect -1577 -1118 -1519 -1106
rect -1319 -130 -1261 -118
rect -1319 -1106 -1307 -130
rect -1273 -1106 -1261 -130
rect -1319 -1118 -1261 -1106
rect -1061 -130 -1003 -118
rect -1061 -1106 -1049 -130
rect -1015 -1106 -1003 -130
rect -1061 -1118 -1003 -1106
rect -803 -130 -745 -118
rect -803 -1106 -791 -130
rect -757 -1106 -745 -130
rect -803 -1118 -745 -1106
rect -545 -130 -487 -118
rect -545 -1106 -533 -130
rect -499 -1106 -487 -130
rect -545 -1118 -487 -1106
rect -287 -130 -229 -118
rect -287 -1106 -275 -130
rect -241 -1106 -229 -130
rect -287 -1118 -229 -1106
rect -29 -130 29 -118
rect -29 -1106 -17 -130
rect 17 -1106 29 -130
rect -29 -1118 29 -1106
rect 229 -130 287 -118
rect 229 -1106 241 -130
rect 275 -1106 287 -130
rect 229 -1118 287 -1106
rect 487 -130 545 -118
rect 487 -1106 499 -130
rect 533 -1106 545 -130
rect 487 -1118 545 -1106
rect 745 -130 803 -118
rect 745 -1106 757 -130
rect 791 -1106 803 -130
rect 745 -1118 803 -1106
rect 1003 -130 1061 -118
rect 1003 -1106 1015 -130
rect 1049 -1106 1061 -130
rect 1003 -1118 1061 -1106
rect 1261 -130 1319 -118
rect 1261 -1106 1273 -130
rect 1307 -1106 1319 -130
rect 1261 -1118 1319 -1106
rect 1519 -130 1577 -118
rect 1519 -1106 1531 -130
rect 1565 -1106 1577 -130
rect 1519 -1118 1577 -1106
rect 1777 -130 1835 -118
rect 1777 -1106 1789 -130
rect 1823 -1106 1835 -130
rect 1777 -1118 1835 -1106
<< mvpdiffc >>
rect -1823 130 -1789 1106
rect -1565 130 -1531 1106
rect -1307 130 -1273 1106
rect -1049 130 -1015 1106
rect -791 130 -757 1106
rect -533 130 -499 1106
rect -275 130 -241 1106
rect -17 130 17 1106
rect 241 130 275 1106
rect 499 130 533 1106
rect 757 130 791 1106
rect 1015 130 1049 1106
rect 1273 130 1307 1106
rect 1531 130 1565 1106
rect 1789 130 1823 1106
rect -1823 -1106 -1789 -130
rect -1565 -1106 -1531 -130
rect -1307 -1106 -1273 -130
rect -1049 -1106 -1015 -130
rect -791 -1106 -757 -130
rect -533 -1106 -499 -130
rect -275 -1106 -241 -130
rect -17 -1106 17 -130
rect 241 -1106 275 -130
rect 499 -1106 533 -130
rect 757 -1106 791 -130
rect 1015 -1106 1049 -130
rect 1273 -1106 1307 -130
rect 1531 -1106 1565 -130
rect 1789 -1106 1823 -130
<< mvnsubdiff >>
rect -1969 1337 1969 1349
rect -1969 1303 -1861 1337
rect 1861 1303 1969 1337
rect -1969 1291 1969 1303
rect -1969 1241 -1911 1291
rect -1969 -1241 -1957 1241
rect -1923 -1241 -1911 1241
rect 1911 1241 1969 1291
rect -1969 -1291 -1911 -1241
rect 1911 -1241 1923 1241
rect 1957 -1241 1969 1241
rect 1911 -1291 1969 -1241
rect -1969 -1303 1969 -1291
rect -1969 -1337 -1861 -1303
rect 1861 -1337 1969 -1303
rect -1969 -1349 1969 -1337
<< mvnsubdiffcont >>
rect -1861 1303 1861 1337
rect -1957 -1241 -1923 1241
rect 1923 -1241 1957 1241
rect -1861 -1337 1861 -1303
<< poly >>
rect -1777 1199 -1577 1215
rect -1777 1165 -1761 1199
rect -1593 1165 -1577 1199
rect -1777 1118 -1577 1165
rect -1519 1199 -1319 1215
rect -1519 1165 -1503 1199
rect -1335 1165 -1319 1199
rect -1519 1118 -1319 1165
rect -1261 1199 -1061 1215
rect -1261 1165 -1245 1199
rect -1077 1165 -1061 1199
rect -1261 1118 -1061 1165
rect -1003 1199 -803 1215
rect -1003 1165 -987 1199
rect -819 1165 -803 1199
rect -1003 1118 -803 1165
rect -745 1199 -545 1215
rect -745 1165 -729 1199
rect -561 1165 -545 1199
rect -745 1118 -545 1165
rect -487 1199 -287 1215
rect -487 1165 -471 1199
rect -303 1165 -287 1199
rect -487 1118 -287 1165
rect -229 1199 -29 1215
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect -229 1118 -29 1165
rect 29 1199 229 1215
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 29 1118 229 1165
rect 287 1199 487 1215
rect 287 1165 303 1199
rect 471 1165 487 1199
rect 287 1118 487 1165
rect 545 1199 745 1215
rect 545 1165 561 1199
rect 729 1165 745 1199
rect 545 1118 745 1165
rect 803 1199 1003 1215
rect 803 1165 819 1199
rect 987 1165 1003 1199
rect 803 1118 1003 1165
rect 1061 1199 1261 1215
rect 1061 1165 1077 1199
rect 1245 1165 1261 1199
rect 1061 1118 1261 1165
rect 1319 1199 1519 1215
rect 1319 1165 1335 1199
rect 1503 1165 1519 1199
rect 1319 1118 1519 1165
rect 1577 1199 1777 1215
rect 1577 1165 1593 1199
rect 1761 1165 1777 1199
rect 1577 1118 1777 1165
rect -1777 71 -1577 118
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 118
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 118
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 118
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 118
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 118
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 118
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 118
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 118
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 118
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -118 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -118 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -118 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -118 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -118 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -118 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -118 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -118 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -118 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -118 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -118 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -118 1777 -71
rect -1777 -1165 -1577 -1118
rect -1777 -1199 -1761 -1165
rect -1593 -1199 -1577 -1165
rect -1777 -1215 -1577 -1199
rect -1519 -1165 -1319 -1118
rect -1519 -1199 -1503 -1165
rect -1335 -1199 -1319 -1165
rect -1519 -1215 -1319 -1199
rect -1261 -1165 -1061 -1118
rect -1261 -1199 -1245 -1165
rect -1077 -1199 -1061 -1165
rect -1261 -1215 -1061 -1199
rect -1003 -1165 -803 -1118
rect -1003 -1199 -987 -1165
rect -819 -1199 -803 -1165
rect -1003 -1215 -803 -1199
rect -745 -1165 -545 -1118
rect -745 -1199 -729 -1165
rect -561 -1199 -545 -1165
rect -745 -1215 -545 -1199
rect -487 -1165 -287 -1118
rect -487 -1199 -471 -1165
rect -303 -1199 -287 -1165
rect -487 -1215 -287 -1199
rect -229 -1165 -29 -1118
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect -229 -1215 -29 -1199
rect 29 -1165 229 -1118
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 29 -1215 229 -1199
rect 287 -1165 487 -1118
rect 287 -1199 303 -1165
rect 471 -1199 487 -1165
rect 287 -1215 487 -1199
rect 545 -1165 745 -1118
rect 545 -1199 561 -1165
rect 729 -1199 745 -1165
rect 545 -1215 745 -1199
rect 803 -1165 1003 -1118
rect 803 -1199 819 -1165
rect 987 -1199 1003 -1165
rect 803 -1215 1003 -1199
rect 1061 -1165 1261 -1118
rect 1061 -1199 1077 -1165
rect 1245 -1199 1261 -1165
rect 1061 -1215 1261 -1199
rect 1319 -1165 1519 -1118
rect 1319 -1199 1335 -1165
rect 1503 -1199 1519 -1165
rect 1319 -1215 1519 -1199
rect 1577 -1165 1777 -1118
rect 1577 -1199 1593 -1165
rect 1761 -1199 1777 -1165
rect 1577 -1215 1777 -1199
<< polycont >>
rect -1761 1165 -1593 1199
rect -1503 1165 -1335 1199
rect -1245 1165 -1077 1199
rect -987 1165 -819 1199
rect -729 1165 -561 1199
rect -471 1165 -303 1199
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect 303 1165 471 1199
rect 561 1165 729 1199
rect 819 1165 987 1199
rect 1077 1165 1245 1199
rect 1335 1165 1503 1199
rect 1593 1165 1761 1199
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect -1761 -1199 -1593 -1165
rect -1503 -1199 -1335 -1165
rect -1245 -1199 -1077 -1165
rect -987 -1199 -819 -1165
rect -729 -1199 -561 -1165
rect -471 -1199 -303 -1165
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
rect 303 -1199 471 -1165
rect 561 -1199 729 -1165
rect 819 -1199 987 -1165
rect 1077 -1199 1245 -1165
rect 1335 -1199 1503 -1165
rect 1593 -1199 1761 -1165
<< locali >>
rect -1957 1303 -1861 1337
rect 1861 1303 1957 1337
rect -1957 1241 -1923 1303
rect 1923 1241 1957 1303
rect -1777 1165 -1761 1199
rect -1593 1165 -1577 1199
rect -1519 1165 -1503 1199
rect -1335 1165 -1319 1199
rect -1261 1165 -1245 1199
rect -1077 1165 -1061 1199
rect -1003 1165 -987 1199
rect -819 1165 -803 1199
rect -745 1165 -729 1199
rect -561 1165 -545 1199
rect -487 1165 -471 1199
rect -303 1165 -287 1199
rect -229 1165 -213 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 213 1165 229 1199
rect 287 1165 303 1199
rect 471 1165 487 1199
rect 545 1165 561 1199
rect 729 1165 745 1199
rect 803 1165 819 1199
rect 987 1165 1003 1199
rect 1061 1165 1077 1199
rect 1245 1165 1261 1199
rect 1319 1165 1335 1199
rect 1503 1165 1519 1199
rect 1577 1165 1593 1199
rect 1761 1165 1777 1199
rect -1823 1106 -1789 1122
rect -1823 114 -1789 130
rect -1565 1106 -1531 1122
rect -1565 114 -1531 130
rect -1307 1106 -1273 1122
rect -1307 114 -1273 130
rect -1049 1106 -1015 1122
rect -1049 114 -1015 130
rect -791 1106 -757 1122
rect -791 114 -757 130
rect -533 1106 -499 1122
rect -533 114 -499 130
rect -275 1106 -241 1122
rect -275 114 -241 130
rect -17 1106 17 1122
rect -17 114 17 130
rect 241 1106 275 1122
rect 241 114 275 130
rect 499 1106 533 1122
rect 499 114 533 130
rect 757 1106 791 1122
rect 757 114 791 130
rect 1015 1106 1049 1122
rect 1015 114 1049 130
rect 1273 1106 1307 1122
rect 1273 114 1307 130
rect 1531 1106 1565 1122
rect 1531 114 1565 130
rect 1789 1106 1823 1122
rect 1789 114 1823 130
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect -1823 -130 -1789 -114
rect -1823 -1122 -1789 -1106
rect -1565 -130 -1531 -114
rect -1565 -1122 -1531 -1106
rect -1307 -130 -1273 -114
rect -1307 -1122 -1273 -1106
rect -1049 -130 -1015 -114
rect -1049 -1122 -1015 -1106
rect -791 -130 -757 -114
rect -791 -1122 -757 -1106
rect -533 -130 -499 -114
rect -533 -1122 -499 -1106
rect -275 -130 -241 -114
rect -275 -1122 -241 -1106
rect -17 -130 17 -114
rect -17 -1122 17 -1106
rect 241 -130 275 -114
rect 241 -1122 275 -1106
rect 499 -130 533 -114
rect 499 -1122 533 -1106
rect 757 -130 791 -114
rect 757 -1122 791 -1106
rect 1015 -130 1049 -114
rect 1015 -1122 1049 -1106
rect 1273 -130 1307 -114
rect 1273 -1122 1307 -1106
rect 1531 -130 1565 -114
rect 1531 -1122 1565 -1106
rect 1789 -130 1823 -114
rect 1789 -1122 1823 -1106
rect -1777 -1199 -1761 -1165
rect -1593 -1199 -1577 -1165
rect -1519 -1199 -1503 -1165
rect -1335 -1199 -1319 -1165
rect -1261 -1199 -1245 -1165
rect -1077 -1199 -1061 -1165
rect -1003 -1199 -987 -1165
rect -819 -1199 -803 -1165
rect -745 -1199 -729 -1165
rect -561 -1199 -545 -1165
rect -487 -1199 -471 -1165
rect -303 -1199 -287 -1165
rect -229 -1199 -213 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 213 -1199 229 -1165
rect 287 -1199 303 -1165
rect 471 -1199 487 -1165
rect 545 -1199 561 -1165
rect 729 -1199 745 -1165
rect 803 -1199 819 -1165
rect 987 -1199 1003 -1165
rect 1061 -1199 1077 -1165
rect 1245 -1199 1261 -1165
rect 1319 -1199 1335 -1165
rect 1503 -1199 1519 -1165
rect 1577 -1199 1593 -1165
rect 1761 -1199 1777 -1165
rect -1957 -1303 -1923 -1241
rect 1923 -1303 1957 -1241
rect -1957 -1337 -1861 -1303
rect 1861 -1337 1957 -1303
<< viali >>
rect -1761 1165 -1593 1199
rect -1503 1165 -1335 1199
rect -1245 1165 -1077 1199
rect -987 1165 -819 1199
rect -729 1165 -561 1199
rect -471 1165 -303 1199
rect -213 1165 -45 1199
rect 45 1165 213 1199
rect 303 1165 471 1199
rect 561 1165 729 1199
rect 819 1165 987 1199
rect 1077 1165 1245 1199
rect 1335 1165 1503 1199
rect 1593 1165 1761 1199
rect -1823 130 -1789 1106
rect -1565 130 -1531 1106
rect -1307 130 -1273 1106
rect -1049 130 -1015 1106
rect -791 130 -757 1106
rect -533 130 -499 1106
rect -275 130 -241 1106
rect -17 130 17 1106
rect 241 130 275 1106
rect 499 130 533 1106
rect 757 130 791 1106
rect 1015 130 1049 1106
rect 1273 130 1307 1106
rect 1531 130 1565 1106
rect 1789 130 1823 1106
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect -1823 -1106 -1789 -130
rect -1565 -1106 -1531 -130
rect -1307 -1106 -1273 -130
rect -1049 -1106 -1015 -130
rect -791 -1106 -757 -130
rect -533 -1106 -499 -130
rect -275 -1106 -241 -130
rect -17 -1106 17 -130
rect 241 -1106 275 -130
rect 499 -1106 533 -130
rect 757 -1106 791 -130
rect 1015 -1106 1049 -130
rect 1273 -1106 1307 -130
rect 1531 -1106 1565 -130
rect 1789 -1106 1823 -130
rect -1761 -1199 -1593 -1165
rect -1503 -1199 -1335 -1165
rect -1245 -1199 -1077 -1165
rect -987 -1199 -819 -1165
rect -729 -1199 -561 -1165
rect -471 -1199 -303 -1165
rect -213 -1199 -45 -1165
rect 45 -1199 213 -1165
rect 303 -1199 471 -1165
rect 561 -1199 729 -1165
rect 819 -1199 987 -1165
rect 1077 -1199 1245 -1165
rect 1335 -1199 1503 -1165
rect 1593 -1199 1761 -1165
<< metal1 >>
rect -1773 1199 -1581 1205
rect -1773 1165 -1761 1199
rect -1593 1165 -1581 1199
rect -1773 1159 -1581 1165
rect -1515 1199 -1323 1205
rect -1515 1165 -1503 1199
rect -1335 1165 -1323 1199
rect -1515 1159 -1323 1165
rect -1257 1199 -1065 1205
rect -1257 1165 -1245 1199
rect -1077 1165 -1065 1199
rect -1257 1159 -1065 1165
rect -999 1199 -807 1205
rect -999 1165 -987 1199
rect -819 1165 -807 1199
rect -999 1159 -807 1165
rect -741 1199 -549 1205
rect -741 1165 -729 1199
rect -561 1165 -549 1199
rect -741 1159 -549 1165
rect -483 1199 -291 1205
rect -483 1165 -471 1199
rect -303 1165 -291 1199
rect -483 1159 -291 1165
rect -225 1199 -33 1205
rect -225 1165 -213 1199
rect -45 1165 -33 1199
rect -225 1159 -33 1165
rect 33 1199 225 1205
rect 33 1165 45 1199
rect 213 1165 225 1199
rect 33 1159 225 1165
rect 291 1199 483 1205
rect 291 1165 303 1199
rect 471 1165 483 1199
rect 291 1159 483 1165
rect 549 1199 741 1205
rect 549 1165 561 1199
rect 729 1165 741 1199
rect 549 1159 741 1165
rect 807 1199 999 1205
rect 807 1165 819 1199
rect 987 1165 999 1199
rect 807 1159 999 1165
rect 1065 1199 1257 1205
rect 1065 1165 1077 1199
rect 1245 1165 1257 1199
rect 1065 1159 1257 1165
rect 1323 1199 1515 1205
rect 1323 1165 1335 1199
rect 1503 1165 1515 1199
rect 1323 1159 1515 1165
rect 1581 1199 1773 1205
rect 1581 1165 1593 1199
rect 1761 1165 1773 1199
rect 1581 1159 1773 1165
rect -1829 1106 -1783 1118
rect -1829 130 -1823 1106
rect -1789 130 -1783 1106
rect -1829 118 -1783 130
rect -1571 1106 -1525 1118
rect -1571 130 -1565 1106
rect -1531 130 -1525 1106
rect -1571 118 -1525 130
rect -1313 1106 -1267 1118
rect -1313 130 -1307 1106
rect -1273 130 -1267 1106
rect -1313 118 -1267 130
rect -1055 1106 -1009 1118
rect -1055 130 -1049 1106
rect -1015 130 -1009 1106
rect -1055 118 -1009 130
rect -797 1106 -751 1118
rect -797 130 -791 1106
rect -757 130 -751 1106
rect -797 118 -751 130
rect -539 1106 -493 1118
rect -539 130 -533 1106
rect -499 130 -493 1106
rect -539 118 -493 130
rect -281 1106 -235 1118
rect -281 130 -275 1106
rect -241 130 -235 1106
rect -281 118 -235 130
rect -23 1106 23 1118
rect -23 130 -17 1106
rect 17 130 23 1106
rect -23 118 23 130
rect 235 1106 281 1118
rect 235 130 241 1106
rect 275 130 281 1106
rect 235 118 281 130
rect 493 1106 539 1118
rect 493 130 499 1106
rect 533 130 539 1106
rect 493 118 539 130
rect 751 1106 797 1118
rect 751 130 757 1106
rect 791 130 797 1106
rect 751 118 797 130
rect 1009 1106 1055 1118
rect 1009 130 1015 1106
rect 1049 130 1055 1106
rect 1009 118 1055 130
rect 1267 1106 1313 1118
rect 1267 130 1273 1106
rect 1307 130 1313 1106
rect 1267 118 1313 130
rect 1525 1106 1571 1118
rect 1525 130 1531 1106
rect 1565 130 1571 1106
rect 1525 118 1571 130
rect 1783 1106 1829 1118
rect 1783 130 1789 1106
rect 1823 130 1829 1106
rect 1783 118 1829 130
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect -1829 -130 -1783 -118
rect -1829 -1106 -1823 -130
rect -1789 -1106 -1783 -130
rect -1829 -1118 -1783 -1106
rect -1571 -130 -1525 -118
rect -1571 -1106 -1565 -130
rect -1531 -1106 -1525 -130
rect -1571 -1118 -1525 -1106
rect -1313 -130 -1267 -118
rect -1313 -1106 -1307 -130
rect -1273 -1106 -1267 -130
rect -1313 -1118 -1267 -1106
rect -1055 -130 -1009 -118
rect -1055 -1106 -1049 -130
rect -1015 -1106 -1009 -130
rect -1055 -1118 -1009 -1106
rect -797 -130 -751 -118
rect -797 -1106 -791 -130
rect -757 -1106 -751 -130
rect -797 -1118 -751 -1106
rect -539 -130 -493 -118
rect -539 -1106 -533 -130
rect -499 -1106 -493 -130
rect -539 -1118 -493 -1106
rect -281 -130 -235 -118
rect -281 -1106 -275 -130
rect -241 -1106 -235 -130
rect -281 -1118 -235 -1106
rect -23 -130 23 -118
rect -23 -1106 -17 -130
rect 17 -1106 23 -130
rect -23 -1118 23 -1106
rect 235 -130 281 -118
rect 235 -1106 241 -130
rect 275 -1106 281 -130
rect 235 -1118 281 -1106
rect 493 -130 539 -118
rect 493 -1106 499 -130
rect 533 -1106 539 -130
rect 493 -1118 539 -1106
rect 751 -130 797 -118
rect 751 -1106 757 -130
rect 791 -1106 797 -130
rect 751 -1118 797 -1106
rect 1009 -130 1055 -118
rect 1009 -1106 1015 -130
rect 1049 -1106 1055 -130
rect 1009 -1118 1055 -1106
rect 1267 -130 1313 -118
rect 1267 -1106 1273 -130
rect 1307 -1106 1313 -130
rect 1267 -1118 1313 -1106
rect 1525 -130 1571 -118
rect 1525 -1106 1531 -130
rect 1565 -1106 1571 -130
rect 1525 -1118 1571 -1106
rect 1783 -130 1829 -118
rect 1783 -1106 1789 -130
rect 1823 -1106 1829 -130
rect 1783 -1118 1829 -1106
rect -1773 -1165 -1581 -1159
rect -1773 -1199 -1761 -1165
rect -1593 -1199 -1581 -1165
rect -1773 -1205 -1581 -1199
rect -1515 -1165 -1323 -1159
rect -1515 -1199 -1503 -1165
rect -1335 -1199 -1323 -1165
rect -1515 -1205 -1323 -1199
rect -1257 -1165 -1065 -1159
rect -1257 -1199 -1245 -1165
rect -1077 -1199 -1065 -1165
rect -1257 -1205 -1065 -1199
rect -999 -1165 -807 -1159
rect -999 -1199 -987 -1165
rect -819 -1199 -807 -1165
rect -999 -1205 -807 -1199
rect -741 -1165 -549 -1159
rect -741 -1199 -729 -1165
rect -561 -1199 -549 -1165
rect -741 -1205 -549 -1199
rect -483 -1165 -291 -1159
rect -483 -1199 -471 -1165
rect -303 -1199 -291 -1165
rect -483 -1205 -291 -1199
rect -225 -1165 -33 -1159
rect -225 -1199 -213 -1165
rect -45 -1199 -33 -1165
rect -225 -1205 -33 -1199
rect 33 -1165 225 -1159
rect 33 -1199 45 -1165
rect 213 -1199 225 -1165
rect 33 -1205 225 -1199
rect 291 -1165 483 -1159
rect 291 -1199 303 -1165
rect 471 -1199 483 -1165
rect 291 -1205 483 -1199
rect 549 -1165 741 -1159
rect 549 -1199 561 -1165
rect 729 -1199 741 -1165
rect 549 -1205 741 -1199
rect 807 -1165 999 -1159
rect 807 -1199 819 -1165
rect 987 -1199 999 -1165
rect 807 -1205 999 -1199
rect 1065 -1165 1257 -1159
rect 1065 -1199 1077 -1165
rect 1245 -1199 1257 -1165
rect 1065 -1205 1257 -1199
rect 1323 -1165 1515 -1159
rect 1323 -1199 1335 -1165
rect 1503 -1199 1515 -1165
rect 1323 -1205 1515 -1199
rect 1581 -1165 1773 -1159
rect 1581 -1199 1593 -1165
rect 1761 -1199 1773 -1165
rect 1581 -1205 1773 -1199
<< properties >>
string FIXED_BBOX -1940 -1320 1940 1320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 2 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1757787870
<< nwell >>
rect -2 -278 804 278
<< pwell >>
rect -2 278 804 550
rect -2 -550 804 -278
<< mvnmos >>
rect 280 364 380 448
rect 580 364 680 448
rect 280 -448 380 -364
rect 580 -448 680 -364
<< mvpmos >>
rect 122 128 222 212
rect 280 128 380 212
rect 438 128 538 212
rect 580 128 680 212
rect 122 -212 222 -128
rect 280 -212 380 -128
rect 438 -212 538 -128
rect 580 -212 680 -128
<< mvndiff >>
rect 222 440 280 448
rect 222 372 234 440
rect 268 372 280 440
rect 222 364 280 372
rect 380 440 580 448
rect 380 372 392 440
rect 568 372 580 440
rect 380 364 580 372
rect 680 440 738 448
rect 680 372 692 440
rect 726 372 738 440
rect 680 364 738 372
rect 222 -372 280 -364
rect 222 -440 234 -372
rect 268 -440 280 -372
rect 222 -448 280 -440
rect 380 -372 580 -364
rect 380 -440 392 -372
rect 568 -440 580 -372
rect 380 -448 580 -440
rect 680 -372 738 -364
rect 680 -440 692 -372
rect 726 -440 738 -372
rect 680 -448 738 -440
<< mvpdiff >>
rect 64 204 122 212
rect 64 136 76 204
rect 110 136 122 204
rect 64 128 122 136
rect 222 204 280 212
rect 222 136 234 204
rect 268 136 280 204
rect 222 128 280 136
rect 380 204 438 212
rect 380 136 392 204
rect 426 136 438 204
rect 380 128 438 136
rect 538 128 580 212
rect 680 204 738 212
rect 680 136 692 204
rect 726 136 738 204
rect 680 128 738 136
rect 64 -136 122 -128
rect 64 -204 76 -136
rect 110 -204 122 -136
rect 64 -212 122 -204
rect 222 -136 280 -128
rect 222 -204 234 -136
rect 268 -204 280 -136
rect 222 -212 280 -204
rect 380 -136 438 -128
rect 380 -204 392 -136
rect 426 -204 438 -136
rect 380 -212 438 -204
rect 538 -212 580 -128
rect 680 -136 738 -128
rect 680 -204 692 -136
rect 726 -204 738 -136
rect 680 -212 738 -204
<< mvndiffc >>
rect 234 372 268 440
rect 392 372 568 440
rect 692 372 726 440
rect 234 -440 268 -372
rect 392 -440 568 -372
rect 692 -440 726 -372
<< mvpdiffc >>
rect 76 136 110 204
rect 234 136 268 204
rect 392 136 426 204
rect 692 136 726 204
rect 76 -204 110 -136
rect 234 -204 268 -136
rect 392 -204 426 -136
rect 692 -204 726 -136
<< mvpsubdiff >>
rect 104 446 142 470
rect 104 412 106 446
rect 140 412 142 446
rect 104 388 142 412
rect 104 -412 142 -388
rect 104 -446 106 -412
rect 140 -446 142 -412
rect 104 -470 142 -446
<< mvnsubdiff >>
rect 64 -66 88 66
rect 504 -66 528 66
<< mvpsubdiffcont >>
rect 106 412 140 446
rect 106 -446 140 -412
<< mvnsubdiffcont >>
rect 88 -66 504 66
<< poly >>
rect 580 520 680 536
rect 580 486 590 520
rect 670 486 680 520
rect 280 448 380 474
rect 580 448 680 486
rect 280 348 380 364
rect 122 307 538 348
rect 580 338 680 364
rect 122 269 318 307
rect 522 269 538 307
rect 122 228 538 269
rect 122 212 222 228
rect 280 212 380 228
rect 438 212 538 228
rect 580 212 680 238
rect 122 102 222 128
rect 280 102 380 128
rect 438 102 538 128
rect 580 80 680 128
rect 580 46 590 80
rect 670 46 680 80
rect 580 30 680 46
rect 580 -46 680 -30
rect 580 -80 590 -46
rect 670 -80 680 -46
rect 122 -128 222 -102
rect 280 -128 380 -102
rect 438 -128 538 -102
rect 580 -128 680 -80
rect 122 -228 222 -212
rect 280 -228 380 -212
rect 438 -228 538 -212
rect 122 -269 538 -228
rect 580 -238 680 -212
rect 122 -307 318 -269
rect 522 -307 538 -269
rect 122 -348 538 -307
rect 280 -364 380 -348
rect 580 -364 680 -338
rect 280 -474 380 -448
rect 580 -486 680 -448
rect 580 -520 590 -486
rect 670 -520 680 -486
rect 580 -536 680 -520
<< polycont >>
rect 590 486 670 520
rect 318 269 522 307
rect 590 46 670 80
rect 590 -80 670 -46
rect 318 -307 522 -269
rect 590 -520 670 -486
<< locali >>
rect 574 486 586 520
rect 234 444 268 456
rect 376 434 392 440
rect 568 434 584 440
rect 376 378 388 434
rect 572 378 584 434
rect 376 372 392 378
rect 568 372 584 378
rect 676 372 692 440
rect 726 372 742 440
rect 76 208 110 220
rect 676 313 742 372
rect 302 307 742 313
rect 302 269 318 307
rect 522 305 742 307
rect 522 271 576 305
rect 684 271 742 305
rect 522 269 742 271
rect 302 263 742 269
rect 234 120 268 132
rect 392 208 426 220
rect 676 204 742 263
rect 676 136 692 204
rect 726 136 742 204
rect 76 66 110 102
rect 392 66 426 102
rect 72 20 88 66
rect 72 -20 82 20
rect 72 -66 88 -20
rect 504 -66 520 66
rect 670 46 686 80
rect 76 -102 110 -66
rect 392 -102 426 -66
rect 574 -80 590 -46
rect 76 -220 110 -208
rect 234 -132 268 -120
rect 392 -220 426 -208
rect 676 -204 692 -136
rect 726 -204 742 -136
rect 676 -263 742 -204
rect 302 -269 742 -263
rect 302 -307 318 -269
rect 522 -271 742 -269
rect 522 -305 576 -271
rect 684 -305 742 -271
rect 522 -307 742 -305
rect 302 -313 742 -307
rect 676 -372 742 -313
rect 376 -378 392 -372
rect 568 -378 584 -372
rect 376 -434 388 -378
rect 572 -434 584 -378
rect 376 -440 392 -434
rect 568 -440 584 -434
rect 676 -440 692 -372
rect 726 -440 742 -372
rect 234 -456 268 -444
rect 574 -520 586 -486
<< viali >>
rect 106 446 140 490
rect 586 486 590 520
rect 590 486 670 520
rect 670 486 692 520
rect 106 412 140 446
rect 106 384 140 412
rect 234 440 268 444
rect 234 372 268 440
rect 388 378 392 434
rect 392 378 568 434
rect 568 378 572 434
rect 76 204 110 208
rect 76 136 110 204
rect 76 102 110 136
rect 234 204 268 372
rect 576 271 684 305
rect 234 136 268 204
rect 234 132 268 136
rect 392 204 426 208
rect 392 136 426 204
rect 392 102 426 136
rect 82 -20 88 20
rect 88 -20 420 20
rect 564 46 590 80
rect 590 46 670 80
rect 76 -136 110 -102
rect 590 -80 670 -46
rect 670 -80 696 -46
rect 76 -204 110 -136
rect 76 -208 110 -204
rect 234 -136 268 -132
rect 234 -204 268 -136
rect 234 -372 268 -204
rect 392 -136 426 -102
rect 392 -204 426 -136
rect 392 -208 426 -204
rect 576 -305 684 -271
rect 106 -412 140 -384
rect 106 -446 140 -412
rect 106 -490 140 -446
rect 234 -440 268 -372
rect 388 -434 392 -378
rect 392 -434 568 -378
rect 568 -434 572 -378
rect 234 -444 268 -440
rect 586 -520 590 -486
rect 590 -520 670 -486
rect 670 -520 692 -486
<< metal1 >>
rect 100 490 480 532
rect 100 384 106 490
rect 140 486 480 490
rect 140 384 146 486
rect 100 372 146 384
rect 228 444 274 456
rect 70 208 116 220
rect 70 102 76 208
rect 110 102 116 208
rect 228 132 234 444
rect 268 132 274 444
rect 376 440 480 486
rect 574 520 704 526
rect 574 486 586 520
rect 692 486 704 520
rect 574 480 704 486
rect 376 434 584 440
rect 376 378 388 434
rect 572 378 584 434
rect 376 372 584 378
rect 564 305 758 311
rect 564 271 576 305
rect 684 271 758 305
rect 564 265 758 271
rect 228 120 274 132
rect 386 208 432 220
rect 70 88 116 102
rect 386 102 392 208
rect 426 102 432 208
rect 386 88 432 102
rect 70 20 432 88
rect 70 -20 82 20
rect 420 -20 432 20
rect 70 -88 432 -20
rect 70 -102 116 -88
rect 70 -208 76 -102
rect 110 -208 116 -102
rect 386 -102 432 -88
rect 70 -220 116 -208
rect 228 -132 274 -120
rect 100 -384 146 -372
rect 100 -490 106 -384
rect 140 -486 146 -384
rect 228 -444 234 -132
rect 268 -444 274 -132
rect 386 -208 392 -102
rect 426 -208 432 -102
rect 386 -220 432 -208
rect 504 80 682 86
rect 504 46 564 80
rect 670 46 682 80
rect 504 40 682 46
rect 504 -265 550 40
rect 710 -40 758 265
rect 578 -46 758 -40
rect 578 -80 590 -46
rect 696 -80 758 -46
rect 578 -86 758 -80
rect 504 -271 696 -265
rect 504 -305 576 -271
rect 684 -305 696 -271
rect 504 -311 696 -305
rect 228 -456 274 -444
rect 376 -378 584 -372
rect 376 -434 388 -378
rect 572 -434 584 -378
rect 376 -440 584 -434
rect 376 -486 480 -440
rect 140 -490 480 -486
rect 100 -532 480 -490
rect 574 -486 704 -480
rect 574 -520 586 -486
rect 692 -520 704 -486
rect 574 -526 704 -520
<< end >>
